module text_difficulty_rom (
    input  logic [8:0] PixelX,
    input  logic [8:0] PixelY,
    output logic [5:0] Data
);

    logic [47:0] data = 48'b00000000000000000000000000000111110000000101010;
    logic [8:0] bitmapIdx;
    logic [1097:0] bitmap;
    logic [2:0] color;

    localparam bit [1097:0] BITMAPS [263] = '{


        // <--- FILE: ASSETS\TEXT\DIFFICULTY\DIFFICULTY.PNG --->

        //tile 0, VRAM 48'b000000000000000000000000000001111100000001010100
        1098'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001,
        1098'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001,
        1098'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001,
        1098'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001,
        1098'b000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000001001001001001001001001001001000000000000010010010010010010010010010010000000000000001000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000001000000000000010010010010010010010010010010000000000000001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000001001001001001000000000000010010010010010010010010010010000000000000001001001001001001000000000000010010010010010010010010010010000000000000001000000000000010010010010010010010010010010000000000000001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000001001001001001,
        1098'b000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000001001001001001000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000001001001001001000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000001001001001001000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000001001001001001000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000001000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000001000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001000000000000000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000001000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001000000000000000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000001000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001000000000000000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000001000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001000000000000000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001001000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001001000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001001000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001001000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000000000000000001001001001001,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000000000000000001001001001001,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000000000000000001001001001001,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000000000000000001001001001001,
        1098'b000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000000000000000001001001001001,
        1098'b000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001,
        1098'b000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001,
        1098'b000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001,
        1098'b000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001,
        1098'b000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000010010010010010010010010010010000000000000000000000000000000010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010000000000000000000000000001001001001001001001001001001,
        1098'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001,
        1098'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001,
        1098'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001,
        1098'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001,
        1098'b001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001,
        1098'b001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001,
        1098'b001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001,
        1098'b001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001,
        1098'b001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000001001001001001000000000010010010010010010010010010010010010010010010010010010010010010000000000001001001001001001001001000000000010010010010010010010010010010010010010010010010010010010010010000000000001001001001000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000001001001001000000000010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000001001001001000000000010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000001001001001000000000010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000001001001001000000000010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000001001001001001000000000010010010010010010010010010000000000001001001001000000000010010010010010010010010010010010010010010010010010010010010010000000000001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000001001001001000000000000010010010010010010010010000000000001001001001001000000000010010010010010010010010010000000000001001001001000000000010010010010010010010010010010010010010010010010010010010010010000000000001001001001000000000000010010010010010010010010000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000001000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000001000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000001000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010010010010010000000000010010010010010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010000000000010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010000000000010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010000000000010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010000000000010010010010010000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010000000000010010010010010000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010000000000010010010010010000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000010010010010010000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000001001001001001000000000010010010010010010010010010000000000001001001001001000000000010010010010010010010010010010010010010010010010010010010010010000000000001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000001001001001000000000000010010010010010010010010010010010010010010010010010010010010000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010010010010010000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010010010010010000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010000000000000000000000000000000000010010010010010010010010010000000000000000000000010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        1098'b001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001
    
    };

    always_comb
    begin
        bitmapIdx = PixelY;
        bitmap    = BITMAPS[bitmapIdx];
        color     = bitmap[3*(365-PixelX) +: 3];
        Data      = data[6*color+0 +: 6];
    end

endmodule
