module text_winner_rom (
    input  logic Tile,
    input  logic [8:0] PixelX,
    input  logic [5:0] PixelY,
    output logic [5:0] Data
);

    logic [48:0] data;
    logic [7:0] bitmapIdx;
    logic [980:0] bitmap;
    logic [2:0] color;

    localparam bit [48:0] DATA [2] = '{


        // <--- FILE: ASSETS\TEXT\WINNER\P1WIN.PNG --->

        //tile 0
        49'b0000000000000000000000001111100000011010100000000,

        // <--- FILE: ASSETS\TEXT\WINNER\P2WIN.PNG --->

        //tile 0
        49'b0000000000000000000000001111100000100000001010101
    
    };

    localparam bit [980:0] BITMAPS [114] = '{


        // <--- FILE: ASSETS\TEXT\WINNER\P1WIN.PNG --->

        //tile 0, VRAM 49'b0000000000000000000000001111100000011010100000000
        981'b000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000,
        981'b000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000,
        981'b000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000,
        981'b000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000,
        981'b000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000,
        981'b000000000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001000001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001000001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001000001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001000001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001000001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001000001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001011011011011011011011001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001011011011011011011011001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001011011011011011011001001001001001001001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001011011011011011011011001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001011011011011011011001001001001001001001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001011011011011011011011001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001011011011011011011001001001001001001001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001011011011011011011011001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001011011011011011011001001001001001001001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001011011011011011011011001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011001001001001001001001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011001001001001001001001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011001001001001001001001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011001001001001001001001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011001001001001001001001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011001001001001001001001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011001001001001001001001001001001001001001001,
        981'b000000000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011001001001001001001001001001001001000000000,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011011011011011011011001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011011011011011011011001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011011011011011011011001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011011011011011011011001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011011011011011011011001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001000000000000000000000000000000000000000000000000001001001001001001011011011011011011011011011011011011011011011011011011001001001001001011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011001001001001001001001001001001001000000000,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001011011011011011011001001001001001001001001001001001000000000,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001011011011011011011001001001001001001001001001001001000000000,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001011011011011011011001001001001001001001001001001001000000000,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001011011011011011011001001001001001001001001001001001000000000,
        981'b000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011001001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011001001001001001001001001001001001001001001001001001001011011011011011011001001001001001001001001001001001000000000,
        981'b000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000,
        981'b000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000,
        981'b000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000,
        981'b000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000,
        981'b000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000,
        981'b000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001000000000,
        981'b000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001000000000,
        981'b000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001000000000,
        981'b000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001000000000,
        981'b000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001000000000,
        981'b000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001000000000,

        // <--- FILE: ASSETS\TEXT\WINNER\P2WIN.PNG --->

        //tile 1, VRAM 49'b0000000000000000000000001111100000100000001010101
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000001000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000001000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000001000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000001000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000001000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000001000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000001000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000010010010010010010010010010010010010000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        981'b001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000,
        981'b001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000,
        981'b001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000,
        981'b001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000,
        981'b001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000,
        981'b001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000
    
    };

    always_comb
    begin
        data      = DATA[Tile];
        bitmapIdx = 7'd57 * data[0] + PixelY;
        bitmap    = BITMAPS[bitmapIdx];
        color     = bitmap[3*(326-PixelX) +: 3];
        Data      = data[6*color+1 +: 6];
    end

endmodule
