module text_title_rom (
    input  logic [8:0] PixelX,
    input  logic [7:0] PixelY,
    output logic [5:0] Data
);

    logic [47:0] data = 48'b00000000000000000000000000000111110101010000000;
    logic [7:0] bitmapIdx;
    logic [1127:0] bitmap;
    logic [2:0] color;

    localparam bit [1127:0] BITMAPS [152] = '{


        // <--- FILE: ASSETS\TEXT\TITLE\TITLE.PNG --->

        //tile 0, VRAM 48'b000000000000000000000000000001111101010100000000
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000000000000000000000001001001001001010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000,
        1128'b000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000,
        1128'b000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000,
        1128'b000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000,
        1128'b000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000,
        1128'b000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000,
        1128'b000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000,
        1128'b000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000,
        1128'b000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000,
        1128'b000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000000000000000000000,
        1128'b000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001000000000000000000000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001001010010010010010010010010010010010010001001001001001001001001001001001001001001001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000,
        1128'b000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000,
        1128'b000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000,
        1128'b000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000,
        1128'b000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000,
        1128'b000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000,
        1128'b000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000,
        1128'b000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001000000000001001001001001001001001001001001001001000000000001001001001001001001001001001001001001001001000000001001001001001001001001001001001001000000000000001001001001001001001001001001001001000000000000000000000000000001001001001001001001001001001001000000000000000001001001001001001001001001001001000000000001001001001001001000000000001001001001001001000001001001001001001001001001001001001001000001001001001001001000001001001001001001000000001001001001001001001000001001001001001001000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001000000000001001001001001001001001001001001001000000000000000000000000000001001001001001001001001001001001000000000001001001001001001001001001001001001001000000000001001001001001001001001001001001000000000001001001001001001001001001001001001001000000000001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010010010010010010010010010010001000000000001010010010010010010010010010010010001000000000001010010010010010010010010010010010010010001000000001010010010010010010010010010010001000000000000001010010010010010010010010010010001000000000000000000000000000001010010010010010010010010010001000000000000000001010010010010010010010010010001000000000001010010010010001000000000001010010010010001001001010010010010010010010010010010010001001001010010010010001001001010010010010001000000001010010010010010001000001010010010010001000000001010010010010010001001010010010010010010010010010010010010010001000000000000000000001010010010010010010010010010010010001000000000001010010010010010010010010010010001000000000000000000000000000001010010010010010010010010010001000000000001010010010010010010010010010010010001000000000001010010010010010010010010010001000000000001010010010010010010010010010010010001000000000001010010010010010010010010010010010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010010010010010010010010010010001001001000001010010010010010010010010010010010001001001000001010010010010010010010010010010010010010001001001001010010010010010010010010010010001001000001001001010010010010010010010010010010001001000000000000000000001001001010010010010010010010010010001001001000001001001010010010010010010010010010001001001000001010010010010001001001001001010010010010001001001010010010010010010010010010010010001001001010010010010001001001010010010010001001001001010010010010010001001001010010010010001001001001010010010010010001001010010010010010010010010010010010010010001001001000000000000001010010010010010010010010010010010001001001001001010010010010010010010010010010001001000000000000000000001001001010010010010010010010010010001001001000001010010010010010010010010010010010001001001001001010010010010010010010010010001001001000001010010010010010010010010010010010001001001000001010010010010010010010010010010010001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001000000000000000000001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001000001010010010010010010001001001010010010010001001001010010010010010010010010010010010001001001010010010010001001001010010010010010010001001010010010010010001001001010010010010001001001001010010010010010001001010010010010010010010010010010010010010001001001000000000000001010010010010010010010010010010010001001001010010010010010010010010010010010010010001000000000000000000001010010010010010010010010010010010010010001000001010010010010010010010010010010010001001001001010010010010010010010010010010010010001000001010010010010010010010010010010010010010001000001010010010010010010010010010010010001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001010010010010010001001001001010010010010001001001010010010010010001001001001010010010010001001001000000000000001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010010010001001001010010010010001001001001001001010010010010001001001001001001001010010010010001001001010010010010010010001001010010010010010001001001010010010010001001001001010010010010010001001010010010010010001001001001001001001001001001001000000000000001001001001001010010010010001001001001001001010010010010010001001001001010010010010001001001000000000000001010010010010001001001001001010010010010001001001001001001010010010010010001001001001001001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001001001001010010010010001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001010010010010010001001001001010010010010001001001010010010010010001001001001010010010010001001001000000000000001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010010010010010001010010010010001001001000000001010010010010001001001001001001001010010010010001001001010010010010010010010001010010010010010001001001010010010010001001001001010010010010010001001010010010010010001001001001001001001001001001001000000000000000000000000001010010010010001001001001001001010010010010010001001001001010010010010001001001000000000000001010010010010001001001001001010010010010001001001000000001010010010010010001001001001001001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001010010010010010001001001001001001001001001001001010010010010010001001001001001001001001001001001000000000000001010010010010001001001001001001001001001001001001010010010010001001001001001010010010010001001001010010010010010010010010001010010010010001001001000000001010010010010001001001001001001001010010010010001001001010010010010010010010001010010010010010001001001010010010010001001001001010010010010010001001010010010010010001001001001001001001001001001001000000000000000000000000001010010010010001001001001001001010010010010010001001001001010010010010001001001000000000000001010010010010001001001001001001001001001001001001000000001010010010010010001001001001001001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010010010001001001001001010010010010001001001010010010010010010010010010010010001001001001001010010010010010010010010010010010001001001001001001010010010010010010010010010010001001001001001001010010010010010010010010010010001001001001000000000000001010010010010001001001001001001001001001001001001010010010010001001001001001010010010010001001001010010010010001010010010010010010010010001001001000000001010010010010001001001000000000001010010010010001001001010010010010001010010010010010010010010001001001010010010010001001001001010010010010010001001010010010010010010010010010010010010001001000000000000000000000000000000001010010010010001001001000000001010010010010010001001001001010010010010001001001000000000000001001001010010010010010010010010010001001001001001000000001010010010010010001001000000000001010010010010001001001001001010010010010001001001010010010010010010010010010010010001001001001001000000001010010010010001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010010010010010010010010010010010010001001001010010010010010010010010010010010010010001001001010010010010010010010010010010010001001001001001001010010010010010010010010010010010001001001001001010010010010010010010010010010010001001001000000000000001010010010010001001001001001001001001001001000001010010010010001001001001001010010010010001001001010010010010001010010010010010010010010001001001000000001010010010010001001001000000000001010010010010001001001010010010010001010010010010010010010010001001001010010010010001001001001010010010010010001001010010010010010010010010010010010010001001000000000000000000000000000000001010010010010001001001000000001010010010010010001001001001010010010010001001001000000000000001001001010010010010010010010010010010010001001001000000001010010010010010001001000000000001010010010010010010010010010010010010010001001001010010010010010010010010010010010010010001001001000000001010010010010001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010010010010010010010010010010001001001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001001001001001001001001001001010010010010001001001001001001001001001001001001010010010010001001001000000000000001010010010010001001001001001001001001001001000001010010010010001001001001001010010010010001001001010010010010001001001010010010010010010001001001000000001010010010010001001001000000000001010010010010001001001010010010010001001001010010010010010010001001001010010010010001001001001010010010010010001001010010010010010001001001001001001001001001000000000000000000000000000000001010010010010001001001000000001010010010010010001001001001010010010010001001001000000000000001001001001001001001001001001010010010010001001001000000001010010010010010001001000000000001010010010010010010010010010010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010010010010010010010010010010001001001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001010010010010010001001001001010010010010001001001010010010010010001001001001010010010010001001001000000000000001010010010010001001001001001010010010010001000001010010010010001001001001001010010010010001001001010010010010001001001010010010010010010001001001000000001010010010010001001001000000000001010010010010001001001010010010010001001001010010010010010010001001001010010010010001001001001010010010010010001001010010010010010001001001001001001001001001000000000000000000000000000000001010010010010001001001000000001010010010010010001001001001010010010010001001001000000000000001010010010010001001001001001010010010010001001001000000001010010010010010001001000000000001010010010010010010010010010010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010010010001001001001001001001001001001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001010010010010010001001001001010010010010001001001010010010010010001001001001010010010010001001001000000000000001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010001001001000000000001010010010010001001001010010010010001001001001010010010010010001001001010010010010001001001001010010010010010001001010010010010010001001001001001001001001001000000000000000000000000000000001010010010010001001001000000001010010010010010001001001001010010010010001001001000000000000001010010010010001001001001001010010010010001001001000000001010010010010010001001000000000001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010010010001001001001001001001001001001000001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001001001010010010010010010010010010010010010001001001010010010010010010010010010010010010010001001001000000000000001010010010010010010010010010010010010010001001001010010010010010010010010010010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010001001001000000000001010010010010001001001010010010010001001001001010010010010010001001001010010010010010010010010010010010010010001001010010010010010010010010010010010010010001000000000000000000000000000000001010010010010001001001000000001010010010010010010010010010010010010010001001001000000000000001010010010010010010010010010010010010010001001001000000001010010010010010001001000000000001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010010010001001001001001001001001001001000001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001001001001010010010010010010010010010010001001001001001001010010010010010010010010010010001001001001000000000000001001001010010010010010010010010010001001001001001001001010010010010010010010010010001001001001001010010010010001001001001001010010010010001001001000000001010010010010001001001000000000001010010010010001001001010010010010001001001001010010010010010001001001001010010010010010010010010010010001001001001010010010010010010010010010010010010010001001001000000000000000000000000001010010010010001001001000000001001001010010010010010010010010010010001001001001000000000000001001001010010010010010010010010010001001001001001000000001010010010010010001001000000000001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000001001001001001001001001000000000001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000001001001001001001001001000000000000001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001000000001001001001001001001001000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000001001001001001001000000001001001001001001001001001001001001001001001001001001001001001001000000000001001001001001001001001001001001000000000000000001001001001001001001001001001001000000000000000000000000000000001001001001001001001001001001001000000000000001001001001001001001001001001001001001000000001001001001001001000000001001001001001001001000000000000001001001001001001000000000000001001001001001001001001001001001001001001000000001001001001001001000000000001001001001001001001001001001001001000000001001001001001001001001001001001001001001001000000000000000000000000000001001001001001001001000000000000000000001001001001001001001001001001001000000000000000000000000000000001001001001001001001001001001001000000000000000000001001001001001001000000000000000001001001001001001000000000001001001001001001001001001001001001001000000001001001001001001001000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000001001001001001001000000001001001001001001001001001001001001001001001001001001001001001001000000000001001001001001001001001001001001000000000000000001001001001001001001001001001001000000000000000000000000000000001001001001001001001001001001001000000000000001001001001001001001001001001001001000000000001001001001001001000000001001001001001001001000000000000001001001001001001000000000000001001001001001001001001001001001001001001000000001001001001001001000000000001001001001001001001001001001001001000000001001001001001001001001001001001001001001001000000000000000000000000000001001001001001001001000000000000000000001001001001001001001001001001001000000000000000000000000000000001001001001001001001001001001001000000000000000000001001001001001001000000000000000001001001001001001000000000001001001001001001000001001001001001001000000001001001001001001001000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1128'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
    
    };

    always_comb
    begin
        bitmapIdx = PixelY;
        bitmap    = BITMAPS[bitmapIdx];
        color     = bitmap[3*(375-PixelX) +: 3];
        Data      = data[6*color+0 +: 6];
    end

endmodule
