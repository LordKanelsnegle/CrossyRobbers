module map_rom (
    input logic [10:0] addr,
    output logic [55:0] data
);

    parameter bit [55:0] ROM [1200] = '{
        //Tile 0 (0,0)
        56'b00000000000000000000000000010000001100001000000100000000,
        //Tile 1 (1,0)
        56'b00000000000000000000000000010000001100001000000100000000,
        //Tile 2 (2,0)
        56'b00000000000000000000000000010000001100001000000100000000,
        //Tile 3 (3,0)
        56'b00000000000000000000000000010000001100001000000100000000,
        //Tile 4 (4,0)
        56'b00000000000000000000000000001100010000001000000100000001,
        //Tile 5 (5,0)
        56'b00000000000000000000100100100000011100011000010100000010,
        //Tile 6 (6,0)
        56'b00000000000000000000000000100100100000010100011000000011,
        //Tile 7 (7,0)
        56'b00000000000000000000000000100100100000010100011000000011,
        //Tile 8 (8,0)
        56'b00000000000000000000100100100000011100010100011000000100,
        //Tile 9 (9,0)
        56'b00000000000000000000001000101000001100000100010000000101,
        //Tile 10 (10,0)
        56'b00000000000000000000001000010000001100000100101000000110,
        //Tile 11 (11,0)
        56'b00000000000000000000001000010000001100000100101000000110,
        //Tile 12 (12,0)
        56'b00000000000000000000001000010000001100000100101000000111,
        //Tile 13 (13,0)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 14 (14,0)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 15 (15,0)
        56'b00000000001000001100110100110000101100010000000100001001,
        //Tile 16 (16,0)
        56'b00000000000000000000000000001000001100000100010000001010,
        //Tile 17 (17,0)
        56'b00000001001001000101000000111100101000010000111000001011,
        //Tile 18 (18,0)
        56'b00000000000000000000000001001100111100111000010000001100,
        //Tile 19 (19,0)
        56'b00000000000000000000000000000001001100111000111100001101,
        //Tile 20 (20,0)
        56'b00000000000000000000000000010000111001001100111100001110,
        //Tile 21 (21,0)
        56'b00000000000000000000000000001000001100000100010000001010,
        //Tile 22 (22,0)
        56'b00000000001000001100000100101100110000110100010000001111,
        //Tile 23 (23,0)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 24 (24,0)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 25 (25,0)
        56'b00000000000000000000100100100000011100011000010100000010,
        //Tile 26 (26,0)
        56'b00000000000000000000000000100100100000010100011000000011,
        //Tile 27 (27,0)
        56'b00000000000000000000000000100100100000010100011000000011,
        //Tile 28 (28,0)
        56'b00000000000000000000000000100100100000010100011000000011,
        //Tile 29 (29,0)
        56'b00000000000000000000000000100100100000010100011000000011,
        //Tile 30 (30,0)
        56'b00000000000000000000100100100000011100010100011000000100,
        //Tile 31 (31,0)
        56'b00000000000000000000000001011101011001010101010000010000,
        //Tile 32 (32,0)
        56'b00000000000000000000000001011101011001010101010000010001,
        //Tile 33 (33,0)
        56'b00000000000000000000000001011101011001010101010000010001,
        //Tile 34 (34,0)
        56'b00000000000000000000000001011101011001010101010000010001,
        //Tile 35 (35,0)
        56'b00000000000000000000000001011101011001010101010000010001,
        //Tile 36 (36,0)
        56'b00000000000000000000000001011101011001010101010000010010,
        //Tile 37 (37,0)
        56'b00000000000000000000000001101101101001100101100000010011,
        //Tile 38 (38,0)
        56'b00000000000000000000000001100001101101101001100100010100,
        //Tile 39 (39,0)
        56'b00000000000000000000000001101101101001100001100100010101,
        //Tile 40 (0,1)
        56'b00000000000000000000000000101000001100000100001000010110,
        //Tile 41 (1,1)
        56'b00000000000000000000000000101000001100000100001000010110,
        //Tile 42 (2,1)
        56'b00000000000000000000000000101000001100000100001000010110,
        //Tile 43 (3,1)
        56'b00000000000000000000000000101000001100000100001000010110,
        //Tile 44 (4,1)
        56'b00000000000000000000000000101000001100000100001000010111,
        //Tile 45 (5,1)
        56'b00000000000000000000000000000001101101100001100100011000,
        //Tile 46 (6,1)
        56'b00000000000000000000000000000001100101101101100000011001,
        //Tile 47 (7,1)
        56'b00000000000000000000000000000001100101101101100000011001,
        //Tile 48 (8,1)
        56'b00000000000000000000000000000001101101100101100000011010,
        //Tile 49 (9,1)
        56'b00000000000000000000000001010101010001011101110000011011,
        //Tile 50 (10,1)
        56'b00000000000000000000000001010101010001110001011100011100,
        //Tile 51 (11,1)
        56'b00000000000000000000000001010101010001110001011100011100,
        //Tile 52 (12,1)
        56'b00000000000000000000000001010101010001110001011100011101,
        //Tile 53 (13,1)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 54 (14,1)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 55 (15,1)
        56'b00000000110000101100110100001100010000001000000100011110,
        //Tile 56 (16,1)
        56'b00000000000000000000000000001000001100000100010000001010,
        //Tile 57 (17,1)
        56'b00000001001001000101000000111100101000010000111000001011,
        //Tile 58 (18,1)
        56'b00000001000001001001000100111101001100010000111000011111,
        //Tile 59 (19,1)
        56'b00000000011100010101110000111100010000111001001100100000,
        //Tile 60 (20,1)
        56'b00000000000001000000111100101000111000010001001100100001,
        //Tile 61 (21,1)
        56'b00000000000000000000000000001000001100000100010000001010,
        //Tile 62 (22,1)
        56'b00000000101100110000001100110100000100010000001000100010,
        //Tile 63 (23,1)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 64 (24,1)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 65 (25,1)
        56'b00000000000000000000000000010100011100100101110100100011,
        //Tile 66 (26,1)
        56'b00000000000000000000000000010100011101110100100100100100,
        //Tile 67 (27,1)
        56'b00000000000000000000000000010100011101110100100100100100,
        //Tile 68 (28,1)
        56'b00000000000000000000000000010100011101110100100100100100,
        //Tile 69 (29,1)
        56'b00000000000000000000000000010100011101110100100100100100,
        //Tile 70 (30,1)
        56'b00000000000000000000000000010100011101110100100100100101,
        //Tile 71 (31,1)
        56'b00000000000000000000101001111000001100000100001000100110,
        //Tile 72 (32,1)
        56'b00000000000000000000101001111000001100000100001000100111,
        //Tile 73 (33,1)
        56'b00000000000000000000000000101000001100000100001000101000,
        //Tile 74 (34,1)
        56'b00000000000000000000000000101000001100000100001000101001,
        //Tile 75 (35,1)
        56'b00000000000000000000101001111000001100000100001000100111,
        //Tile 76 (36,1)
        56'b00000000000000000000101001111000001100000100001000101010,
        //Tile 77 (37,1)
        56'b00000000000000000000000000000001101101100001100100011000,
        //Tile 78 (38,1)
        56'b00000000001100010000111000000100111100101000001000101011,
        //Tile 79 (39,1)
        56'b00000000000000000000000000000001101101100101100000011010,
        //Tile 80 (0,2)
        56'b00000000000000000000101001111000001100000100001000101100,
        //Tile 81 (1,2)
        56'b00000000000000000000000000010000000100001001111000101101,
        //Tile 82 (2,2)
        56'b00000000000000000000000000010000000100001001111000101110,
        //Tile 83 (3,2)
        56'b00000000000000000000101001111000001100000100001000101111,
        //Tile 84 (4,2)
        56'b00000000000000000000101001111000001100000100001000110000,
        //Tile 85 (5,2)
        56'b00000000000000010000111000000100111100101000001000110001,
        //Tile 86 (6,2)
        56'b00000000000000010000000100111000101000111100001000110010,
        //Tile 87 (7,2)
        56'b00000000000000000001100001010001011001011101010100110011,
        //Tile 88 (8,2)
        56'b00101100110000101000100001100001100100010000001000110100,
        //Tile 89 (9,2)
        56'b00000000000000000000000001010101010001011101110000110101,
        //Tile 90 (10,2)
        56'b00000000000000000000000000001000001100000100101000110110,
        //Tile 91 (11,2)
        56'b00000000000000000000000000001000001100000100101000110110,
        //Tile 92 (12,2)
        56'b00000000000000000000000001010101010001011101110000110101,
        //Tile 93 (13,2)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 94 (14,2)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 95 (15,2)
        56'b00000000001000001100110100110000101100010000000100001001,
        //Tile 96 (16,2)
        56'b00000000000000000000000000001000001100000100010000110111,
        //Tile 97 (17,2)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 98 (18,2)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 99 (19,2)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 100 (20,2)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 101 (21,2)
        56'b00000000000000000000000000001000010000000100001100111001,
        //Tile 102 (22,2)
        56'b00000000001000001100000100101100110000110100010000001111,
        //Tile 103 (23,2)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 104 (24,2)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 105 (25,2)
        56'b01011001111100100101101000011101110100010000001000111010,
        //Tile 106 (26,2)
        56'b01100001101101100100111000010000111100101000001000111011,
        //Tile 107 (27,2)
        56'b01100001101101100100010000111000101000111100001000111100,
        //Tile 108 (28,2)
        56'b00000001111000010000111000000100111100101000001000111101,
        //Tile 109 (29,2)
        56'b00000001111000010000000100111000101000111100001000111110,
        //Tile 110 (30,2)
        56'b00000000111001011101000001110100011100010000001000111111,
        //Tile 111 (31,2)
        56'b00000000000000000000101001111000001100000100001000100110,
        //Tile 112 (32,2)
        56'b00000000000000000000101001111000001100000100001000101010,
        //Tile 113 (33,2)
        56'b00000000000000000000000000010000000100001001111000101101,
        //Tile 114 (34,2)
        56'b00000000000000000000000000010000000100001001111000101110,
        //Tile 115 (35,2)
        56'b00000000000000000000101001111000001100000100001000100110,
        //Tile 116 (36,2)
        56'b00000000000000000000101001111000001100000100001000101010,
        //Tile 117 (37,2)
        56'b01100001101101100100111000010000111100101000001001000000,
        //Tile 118 (38,2)
        56'b00000100101001000100110101100101100000010000001001000001,
        //Tile 119 (39,2)
        56'b00000000001100010000111000000100111100101000001000101011,
        //Tile 120 (0,3)
        56'b00000000000000000000000000000000001100001000000101000010,
        //Tile 121 (1,3)
        56'b00000000000000000000000000000100010000001001111001000011,
        //Tile 122 (2,3)
        56'b00000000000000000000000000000100001000010001111001000100,
        //Tile 123 (3,3)
        56'b00000000000000000000000000000000001100000100001001000101,
        //Tile 124 (4,3)
        56'b00000000000000000000000000000000001100001000000101000010,
        //Tile 125 (5,3)
        56'b00000000000000000000000000000001101101100001100100011000,
        //Tile 126 (6,3)
        56'b00000000000000000000000000000001101101100101100000011010,
        //Tile 127 (7,3)
        56'b00000001101001010001000001100001011001011101010101000110,
        //Tile 128 (8,3)
        56'b00000000000000000000000000000001101101100001100101000111,
        //Tile 129 (9,3)
        56'b00000000000000000000000001010101010001011101110000110101,
        //Tile 130 (10,3)
        56'b00000000000000000000000000001000001100000100101000110110,
        //Tile 131 (11,3)
        56'b00000000000000000000000000001000001100000100101000110110,
        //Tile 132 (12,3)
        56'b00000000000000000000000001010101010001011101110000110101,
        //Tile 133 (13,3)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 134 (14,3)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 135 (15,3)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 136 (16,3)
        56'b00000000110000001100101100110100000100010000001001001000,
        //Tile 137 (17,3)
        56'b00000000001100110000101100000100110100001000010001001001,
        //Tile 138 (18,3)
        56'b00000000111001001100111100001100010000001000000101001010,
        //Tile 139 (19,3)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 140 (20,3)
        56'b00000000110000001100101100110100000100010000001001001000,
        //Tile 141 (21,3)
        56'b00000000001100110000101100000100110100001000010001001001,
        //Tile 142 (22,3)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 143 (23,3)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 144 (24,3)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 145 (25,3)
        56'b00000000000000000000000000010100011100100101110101001011,
        //Tile 146 (26,3)
        56'b00000000000000000000000000000001100001101101100101001100,
        //Tile 147 (27,3)
        56'b00000000000000000000000000000001100001101101100101001101,
        //Tile 148 (28,3)
        56'b00000000000000000000000000010100011100100101110100100011,
        //Tile 149 (29,3)
        56'b00000000000000000000000000010100011101110100100100100100,
        //Tile 150 (30,3)
        56'b00000000000000000000000000010100011101110100100100100101,
        //Tile 151 (31,3)
        56'b00000000000000000000000000000000001100000100001001000101,
        //Tile 152 (32,3)
        56'b00000000000000000000000000000000001100001000000101000010,
        //Tile 153 (33,3)
        56'b00000000000000000000000000000100010000001001111001000011,
        //Tile 154 (34,3)
        56'b00000000000000000000000000000100001000010001111001000100,
        //Tile 155 (35,3)
        56'b00000000000000000000000000000000001100000100001001000101,
        //Tile 156 (36,3)
        56'b00000000000000000000000000000000001100001000000101000010,
        //Tile 157 (37,3)
        56'b00000000000000000000000000000001100001101101100101001100,
        //Tile 158 (38,3)
        56'b00000000000000000000000000000001100101101101100000011001,
        //Tile 159 (39,3)
        56'b00000000000000000000000000000001101101100101100000011010,
        //Tile 160 (0,4)
        56'b00111000001100111101001110000000010000001000000101001110,
        //Tile 161 (1,4)
        56'b00000000000000000000000000001000001100000100010001001111,
        //Tile 162 (2,4)
        56'b00000000000000000000000000001000010000000100001101010000,
        //Tile 163 (3,4)
        56'b00000000110000001100101100110100000100010000001001001000,
        //Tile 164 (4,4)
        56'b00000000001100110000101100000100110100001000010001001001,
        //Tile 165 (5,4)
        56'b00111000001100111101001110000000010000001000000101001110,
        //Tile 166 (6,4)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 167 (7,4)
        56'b00000000000000000000000000001000001100000100010001010001,
        //Tile 168 (8,4)
        56'b00000000111001001100111100001100010000001000000101001010,
        //Tile 169 (9,4)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 170 (10,4)
        56'b00000000000000000000000000001000001100000100010001010010,
        //Tile 171 (11,4)
        56'b00000000000000000000000000001000010000000100001101010011,
        //Tile 172 (12,4)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 173 (13,4)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 174 (14,4)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 175 (15,4)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 176 (16,4)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 177 (17,4)
        56'b00000000000010001110001010000100001100001000000101010100,
        //Tile 178 (18,4)
        56'b00000000000010001010010000000010001110000100000101010101,
        //Tile 179 (19,4)
        56'b00000000000000000000000000000000000010001110000101010110,
        //Tile 180 (20,4)
        56'b00000000000000000000000000000010001100000110000101010111,
        //Tile 181 (21,4)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 182 (22,4)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 183 (23,4)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 184 (24,4)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 185 (25,4)
        56'b00111000001100111101001110000000010000001000000101001110,
        //Tile 186 (26,4)
        56'b00000000000000000000000000001000001100000100010001001111,
        //Tile 187 (27,4)
        56'b00000000000000000000000000001000010000000100001101010000,
        //Tile 188 (28,4)
        56'b00111000001100111101001110000000010000001000000101001110,
        //Tile 189 (29,4)
        56'b00000000110000001100101100110100000100010000001001001000,
        //Tile 190 (30,4)
        56'b00000000001100110000101100000100110100001000010001001001,
        //Tile 191 (31,4)
        56'b00111000001100111101001110000000010000001000000101001110,
        //Tile 192 (32,4)
        56'b00111000111100001101000000101000010000001000000101011000,
        //Tile 193 (33,4)
        56'b00000000000000000000000000001000001100000100010001001111,
        //Tile 194 (34,4)
        56'b00000000000000000000000000001000010000000100001101010000,
        //Tile 195 (35,4)
        56'b00111000111100001101000000101000010000001000000101011000,
        //Tile 196 (36,4)
        56'b00111000001100111101001110000000010000001000000101001110,
        //Tile 197 (37,4)
        56'b00000000000000000000000000001000001100000100010001010001,
        //Tile 198 (38,4)
        56'b00000000110000001100101100110100000100010000001001001000,
        //Tile 199 (39,4)
        56'b00000000001100110000101100000100110100001000010001001001,
        //Tile 200 (0,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 201 (1,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 202 (2,5)
        56'b00000000000000000000000000010000001100001000000101011001,
        //Tile 203 (3,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 204 (4,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 205 (5,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 206 (6,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 207 (7,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 208 (8,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 209 (9,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 210 (10,5)
        56'b00000000000000000000000000001000001100000100010001010010,
        //Tile 211 (11,5)
        56'b00000000000000000000000000001000010000000100001101010011,
        //Tile 212 (12,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 213 (13,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 214 (14,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 215 (15,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 216 (16,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 217 (17,5)
        56'b00001000010000001100000110001000000010001110000101011010,
        //Tile 218 (18,5)
        56'b00000000010010010100000010000110001110001010010001011011,
        //Tile 219 (19,5)
        56'b00000000000000010000001010000100000010001010001101011100,
        //Tile 220 (20,5)
        56'b00000000000000001000010000001100000010000110001101011101,
        //Tile 221 (21,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 222 (22,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 223 (23,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 224 (24,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 225 (25,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 226 (26,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 227 (27,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 228 (28,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 229 (29,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 230 (30,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 231 (31,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 232 (32,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 233 (33,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 234 (34,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 235 (35,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 236 (36,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 237 (37,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 238 (38,5)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 239 (39,5)
        56'b00000000000000000000000000010000001100001000000101011001,
        //Tile 240 (0,6)
        56'b00000001111101000001101000001100010000001000000101011110,
        //Tile 241 (1,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 242 (2,6)
        56'b00000000000000000000000000001100010000001000000101011111,
        //Tile 243 (3,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 244 (4,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 245 (5,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 246 (6,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 247 (7,6)
        56'b00000001111101000001101000001100010000001000000101011110,
        //Tile 248 (8,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 249 (9,6)
        56'b00000000000000000000000000010000001100001000000101100000,
        //Tile 250 (10,6)
        56'b00000000000000000000000000001000001100000100010001010010,
        //Tile 251 (11,6)
        56'b00000000000000000000000000001000010000000100001101010011,
        //Tile 252 (12,6)
        56'b00000000000000000000000000010000001100001000000101100000,
        //Tile 253 (13,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 254 (14,6)
        56'b00000001111101000001101000001100010000001000000101011110,
        //Tile 255 (15,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 256 (16,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 257 (17,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 258 (18,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 259 (19,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 260 (20,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 261 (21,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 262 (22,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 263 (23,6)
        56'b00000001111101000001101000001100010000001000000101100001,
        //Tile 264 (24,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 265 (25,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 266 (26,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 267 (27,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 268 (28,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 269 (29,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 270 (30,6)
        56'b00000001111101000001101000001100010000001000000101100001,
        //Tile 271 (31,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 272 (32,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 273 (33,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 274 (34,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 275 (35,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 276 (36,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 277 (37,6)
        56'b00000001111101000001101000001100010000001000000101100001,
        //Tile 278 (38,6)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 279 (39,6)
        56'b00000000000000000000000000001100010000001000000101011111,
        //Tile 280 (0,7)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 281 (1,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 282 (2,7)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 283 (3,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 284 (4,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 285 (5,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 286 (6,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 287 (7,7)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 288 (8,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 289 (9,7)
        56'b00000000000000000000000000010000001100001000000101100011,
        //Tile 290 (10,7)
        56'b00000000000000000000000000001000001100000100010001010010,
        //Tile 291 (11,7)
        56'b00000000000000000000000000001000010000000100001101010011,
        //Tile 292 (12,7)
        56'b00000000000000000000000000010000001100001000000101100011,
        //Tile 293 (13,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 294 (14,7)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 295 (15,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 296 (16,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 297 (17,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 298 (18,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 299 (19,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 300 (20,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 301 (21,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 302 (22,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 303 (23,7)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 304 (24,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 305 (25,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 306 (26,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 307 (27,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 308 (28,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 309 (29,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 310 (30,7)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 311 (31,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 312 (32,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 313 (33,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 314 (34,7)
        56'b00010001011100101001011000001101010100001000000101100100,
        //Tile 315 (35,7)
        56'b00000000000000000001100000001101100100001000000101100101,
        //Tile 316 (36,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 317 (37,7)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 318 (38,7)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 319 (39,7)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 320 (0,8)
        56'b00000000000000000000000000001000000100001100010001100110,
        //Tile 321 (1,8)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 322 (2,8)
        56'b00000000000000000000000000001000000100001100010001100110,
        //Tile 323 (3,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 324 (4,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 325 (5,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 326 (6,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 327 (7,8)
        56'b00000000000000000000000000001000000100001100010001100111,
        //Tile 328 (8,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 329 (9,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 330 (10,8)
        56'b00000000000000000000000000001000001100000100010001001111,
        //Tile 331 (11,8)
        56'b00000000000000000000000000001000010000000100001101010000,
        //Tile 332 (12,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 333 (13,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 334 (14,8)
        56'b00000000000000000000000000001000000100001100010001100111,
        //Tile 335 (15,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 336 (16,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 337 (17,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 338 (18,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 339 (19,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 340 (20,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 341 (21,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 342 (22,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 343 (23,8)
        56'b00000000000000000000000000001000000100001100010001101000,
        //Tile 344 (24,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 345 (25,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 346 (26,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 347 (27,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 348 (28,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 349 (29,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 350 (30,8)
        56'b00000000000000000000000000001000000100001100010001101000,
        //Tile 351 (31,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 352 (32,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 353 (33,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 354 (34,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 355 (35,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 356 (36,8)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 357 (37,8)
        56'b00000000000000000000000000001000000100001100010001101001,
        //Tile 358 (38,8)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 359 (39,8)
        56'b00000000000000000000000000001000000100001100010001101010,
        //Tile 360 (0,9)
        56'b00000000000000000000000000001000001100000100010001101011,
        //Tile 361 (1,9)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 362 (2,9)
        56'b00000000000000000000000000001000000100001100010001101100,
        //Tile 363 (3,9)
        56'b00000000000000000000000000000000101000001000010001101101,
        //Tile 364 (4,9)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 365 (5,9)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 366 (6,9)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 367 (7,9)
        56'b00000000000000000000000000000000101000010000001001110000,
        //Tile 368 (8,9)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 369 (9,9)
        56'b00000000000000000000000000000000000000101000001001110001,
        //Tile 370 (10,9)
        56'b00000000000000000000000000000000000000101000001001110001,
        //Tile 371 (11,9)
        56'b00000000000000000000000000000000000000101000001001110001,
        //Tile 372 (12,9)
        56'b00000000000000000000000000000000000000101000001001110001,
        //Tile 373 (13,9)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 374 (14,9)
        56'b00000000000000000000000000000000101000010000001001110010,
        //Tile 375 (15,9)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 376 (16,9)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 377 (17,9)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 378 (18,9)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 379 (19,9)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 380 (20,9)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 381 (21,9)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 382 (22,9)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 383 (23,9)
        56'b00000000000000000000000000000000101000010000001001110011,
        //Tile 384 (24,9)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 385 (25,9)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 386 (26,9)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 387 (27,9)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 388 (28,9)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 389 (29,9)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 390 (30,9)
        56'b00000000000000000000000000000000101000010000001001110100,
        //Tile 391 (31,9)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 392 (32,9)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 393 (33,9)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 394 (34,9)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 395 (35,9)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 396 (36,9)
        56'b00000000000000000000000000000000000000101000001001110101,
        //Tile 397 (37,9)
        56'b00000000000000000000000000001000001100000100010001110110,
        //Tile 398 (38,9)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 399 (39,9)
        56'b00000000000000000000000000001000000100001100010001101100,
        //Tile 400 (0,10)
        56'b00000000000000000000000000000000000000101000001001110111,
        //Tile 401 (1,10)
        56'b00000000000000000000000000000000000000001000101001111000,
        //Tile 402 (2,10)
        56'b00000000000000000000000000000000101000010000001001111001,
        //Tile 403 (3,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 404 (4,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 405 (5,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 406 (6,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 407 (7,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 408 (8,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 409 (9,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 410 (10,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 411 (11,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 412 (12,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 413 (13,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 414 (14,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 415 (15,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 416 (16,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 417 (17,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 418 (18,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 419 (19,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 420 (20,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 421 (21,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 422 (22,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 423 (23,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 424 (24,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 425 (25,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 426 (26,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 427 (27,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 428 (28,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 429 (29,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 430 (30,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 431 (31,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 432 (32,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 433 (33,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 434 (34,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 435 (35,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 436 (36,10)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 437 (37,10)
        56'b00000000000000000000000000000000000000101000001001110111,
        //Tile 438 (38,10)
        56'b00000000000000000000000000000000000000001000101001111000,
        //Tile 439 (39,10)
        56'b00000000000000000000000000000000101000010000001001111001,
        //Tile 440 (0,11)
        56'b00000000000000000000000000000001000000101000001001111011,
        //Tile 441 (1,11)
        56'b00000000000000000000000000000000000000001000101001111000,
        //Tile 442 (2,11)
        56'b00000000000000000000000000000001000000101000001001111100,
        //Tile 443 (3,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 444 (4,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 445 (5,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 446 (6,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 447 (7,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 448 (8,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 449 (9,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 450 (10,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 451 (11,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 452 (12,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 453 (13,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 454 (14,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 455 (15,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 456 (16,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 457 (17,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 458 (18,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 459 (19,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 460 (20,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 461 (21,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 462 (22,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 463 (23,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 464 (24,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 465 (25,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 466 (26,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 467 (27,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 468 (28,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 469 (29,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 470 (30,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 471 (31,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 472 (32,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 473 (33,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 474 (34,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 475 (35,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 476 (36,11)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 477 (37,11)
        56'b00000000000000000000000000000001000000101000001001111011,
        //Tile 478 (38,11)
        56'b00000000000000000000000000000000000000001000101001111000,
        //Tile 479 (39,11)
        56'b00000000000000000000000000000001000000101000001001111100,
        //Tile 480 (0,12)
        56'b00000000000000000000000000000001000000101000001001111110,
        //Tile 481 (1,12)
        56'b00000000000000000000000000000000000000001000101001111000,
        //Tile 482 (2,12)
        56'b00000000000000000000000000000001000000101000001001111111,
        //Tile 483 (3,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 484 (4,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 485 (5,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 486 (6,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 487 (7,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 488 (8,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 489 (9,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 490 (10,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 491 (11,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 492 (12,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 493 (13,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 494 (14,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 495 (15,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 496 (16,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 497 (17,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 498 (18,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 499 (19,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 500 (20,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 501 (21,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 502 (22,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 503 (23,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 504 (24,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 505 (25,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 506 (26,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 507 (27,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 508 (28,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 509 (29,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 510 (30,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 511 (31,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 512 (32,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 513 (33,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 514 (34,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 515 (35,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 516 (36,12)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 517 (37,12)
        56'b00000000000000000000000000000001000000101000001001111110,
        //Tile 518 (38,12)
        56'b00000000000000000000000000000000000000001000101001111000,
        //Tile 519 (39,12)
        56'b00000000000000000000000000000001000000101000001001111111,
        //Tile 520 (0,13)
        56'b00000000000000000000000000000000000000101000001010000001,
        //Tile 521 (1,13)
        56'b00000000000000000000000000000000000000101000001010000010,
        //Tile 522 (2,13)
        56'b00000000000000000000000000000000000000101000001010000011,
        //Tile 523 (3,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 524 (4,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 525 (5,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 526 (6,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 527 (7,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 528 (8,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 529 (9,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 530 (10,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 531 (11,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 532 (12,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 533 (13,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 534 (14,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 535 (15,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 536 (16,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 537 (17,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 538 (18,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 539 (19,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 540 (20,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 541 (21,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 542 (22,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 543 (23,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 544 (24,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 545 (25,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 546 (26,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 547 (27,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 548 (28,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 549 (29,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 550 (30,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 551 (31,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 552 (32,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 553 (33,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 554 (34,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 555 (35,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 556 (36,13)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 557 (37,13)
        56'b00000000000000000000000000000000000000101000001010000001,
        //Tile 558 (38,13)
        56'b00000000000000000000000000000000000000101000001010000010,
        //Tile 559 (39,13)
        56'b00000000000000000000000000000000000000101000001010000011,
        //Tile 560 (0,14)
        56'b00000000000000000000000000001100000100010000001010000100,
        //Tile 561 (1,14)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 562 (2,14)
        56'b00000000000000000000000000001100000100001000010010000101,
        //Tile 563 (3,14)
        56'b00000000000000000000000000000000000000101000001010000110,
        //Tile 564 (4,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 565 (5,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 566 (6,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 567 (7,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 568 (8,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 569 (9,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 570 (10,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 571 (11,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 572 (12,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 573 (13,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 574 (14,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 575 (15,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 576 (16,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 577 (17,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 578 (18,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 579 (19,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 580 (20,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 581 (21,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 582 (22,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 583 (23,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 584 (24,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 585 (25,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 586 (26,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 587 (27,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 588 (28,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 589 (29,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 590 (30,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 591 (31,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 592 (32,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 593 (33,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 594 (34,14)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 595 (35,14)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 596 (36,14)
        56'b00000000000000000000000000000000000000101000001010001001,
        //Tile 597 (37,14)
        56'b00000000000000000000000000001100000100010000001010000100,
        //Tile 598 (38,14)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 599 (39,14)
        56'b00000000000000000000000000001100000100001000010010000101,
        //Tile 600 (0,15)
        56'b00000000000000000000000000001000001100000100010010001010,
        //Tile 601 (1,15)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 602 (2,15)
        56'b00000000000000000000000000001000001100000100010010001011,
        //Tile 603 (3,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 604 (4,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 605 (5,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 606 (6,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 607 (7,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 608 (8,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 609 (9,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 610 (10,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 611 (11,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 612 (12,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 613 (13,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 614 (14,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 615 (15,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 616 (16,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 617 (17,15)
        56'b00000000000000000000000000001000001100000100010010001100,
        //Tile 618 (18,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 619 (19,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 620 (20,15)
        56'b00000000000000000000000000001000001100000100010010001100,
        //Tile 621 (21,15)
        56'b00000000000000000000000000001000001100000100010010001101,
        //Tile 622 (22,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 623 (23,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 624 (24,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 625 (25,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 626 (26,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 627 (27,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 628 (28,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 629 (29,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 630 (30,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 631 (31,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 632 (32,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 633 (33,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 634 (34,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 635 (35,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 636 (36,15)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 637 (37,15)
        56'b00000000000000000000000000001100000100010000001010001110,
        //Tile 638 (38,15)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 639 (39,15)
        56'b00000000000000000000000000001100000100010000001010001111,
        //Tile 640 (0,16)
        56'b00000001111101000001101000001100010000001000000101011110,
        //Tile 641 (1,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 642 (2,16)
        56'b00000000000000000000000000001100010000001000000101011111,
        //Tile 643 (3,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 644 (4,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 645 (5,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 646 (6,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 647 (7,16)
        56'b00000001111101000001101000001100010000001000000101011110,
        //Tile 648 (8,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 649 (9,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 650 (10,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 651 (11,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 652 (12,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 653 (13,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 654 (14,16)
        56'b00000001111101000001101000001100010000001000000101011110,
        //Tile 655 (15,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 656 (16,16)
        56'b00111000001100111101001110000000010000001000000101001110,
        //Tile 657 (17,16)
        56'b00000000110000001100101100001000110100000100010010010000,
        //Tile 658 (18,16)
        56'b00000000001100110000101100001000000100010000110110010001,
        //Tile 659 (19,16)
        56'b00000000110000001100101100001000110100000100010010010000,
        //Tile 660 (20,16)
        56'b00000000001100110000101100001000000100010000110110010001,
        //Tile 661 (21,16)
        56'b00111000001100111101001110000000010000001000000101001110,
        //Tile 662 (22,16)
        56'b00000000111001001100111100001100010000001000000101001010,
        //Tile 663 (23,16)
        56'b00000001111101000001101000001100010000001000000101011110,
        //Tile 664 (24,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 665 (25,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 666 (26,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 667 (27,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 668 (28,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 669 (29,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 670 (30,16)
        56'b00000001111101000001101000001100010000001000000101100001,
        //Tile 671 (31,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 672 (32,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 673 (33,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 674 (34,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 675 (35,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 676 (36,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 677 (37,16)
        56'b00000001111101000001101000001100010000001000000101100001,
        //Tile 678 (38,16)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 679 (39,16)
        56'b00000000000000000000000000001100010000001000000101011111,
        //Tile 680 (0,17)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 681 (1,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 682 (2,17)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 683 (3,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 684 (4,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 685 (5,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 686 (6,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 687 (7,17)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 688 (8,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 689 (9,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 690 (10,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 691 (11,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 692 (12,17)
        56'b00000000000000000001100000001101100100001000000101100101,
        //Tile 693 (13,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 694 (14,17)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 695 (15,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 696 (16,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 697 (17,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 698 (18,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 699 (19,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 700 (20,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 701 (21,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 702 (22,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 703 (23,17)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 704 (24,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 705 (25,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 706 (26,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 707 (27,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 708 (28,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 709 (29,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 710 (30,17)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 711 (31,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 712 (32,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 713 (33,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 714 (34,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 715 (35,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 716 (36,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 717 (37,17)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 718 (38,17)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 719 (39,17)
        56'b00000000000000000000000000001100010000001000000101100010,
        //Tile 720 (0,18)
        56'b00000000000000000000000000001000000100001100010001100110,
        //Tile 721 (1,18)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 722 (2,18)
        56'b00000000000000000000000000001000000100001100010001100110,
        //Tile 723 (3,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 724 (4,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 725 (5,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 726 (6,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 727 (7,18)
        56'b00000000000000000000000000001000000100001100010001100111,
        //Tile 728 (8,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 729 (9,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 730 (10,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 731 (11,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 732 (12,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 733 (13,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 734 (14,18)
        56'b00000000000000000000000000001000000100001100010001100111,
        //Tile 735 (15,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 736 (16,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 737 (17,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 738 (18,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 739 (19,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 740 (20,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 741 (21,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 742 (22,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 743 (23,18)
        56'b00000000000000000000000000001000000100001100010001100111,
        //Tile 744 (24,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 745 (25,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 746 (26,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 747 (27,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 748 (28,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 749 (29,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 750 (30,18)
        56'b00000000000000000000000000001000000100001100010001101000,
        //Tile 751 (31,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 752 (32,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 753 (33,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 754 (34,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 755 (35,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 756 (36,18)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 757 (37,18)
        56'b00000000000000000000000000001000000100001100010001101001,
        //Tile 758 (38,18)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 759 (39,18)
        56'b00000000000000000000000000001000000100001100010001101010,
        //Tile 760 (0,19)
        56'b00000000000000000000000000001000001100000100010001101011,
        //Tile 761 (1,19)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 762 (2,19)
        56'b00000000000000000000000000001000000100001100010001101100,
        //Tile 763 (3,19)
        56'b00000000000000000000000000000000101000001000010001101101,
        //Tile 764 (4,19)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 765 (5,19)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 766 (6,19)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 767 (7,19)
        56'b00000000000000000000000000000000101000010000001001110000,
        //Tile 768 (8,19)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 769 (9,19)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 770 (10,19)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 771 (11,19)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 772 (12,19)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 773 (13,19)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 774 (14,19)
        56'b00000000000000000000000000000000101000010000001001110010,
        //Tile 775 (15,19)
        56'b00000000000000010001011101011001010100101000001010010010,
        //Tile 776 (16,19)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 777 (17,19)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 778 (18,19)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 779 (19,19)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 780 (20,19)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 781 (21,19)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 782 (22,19)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 783 (23,19)
        56'b00000000000000000000000000000000101000010000001001110000,
        //Tile 784 (24,19)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 785 (25,19)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 786 (26,19)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 787 (27,19)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 788 (28,19)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 789 (29,19)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 790 (30,19)
        56'b00000000000000000000000000000000101000010000001001110100,
        //Tile 791 (31,19)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 792 (32,19)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 793 (33,19)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 794 (34,19)
        56'b00000000000000000000000000000000000000101000001001101110,
        //Tile 795 (35,19)
        56'b00000000000000000000000000000000000000101000001001101111,
        //Tile 796 (36,19)
        56'b00000000000000000000000000000000000000101000001001110101,
        //Tile 797 (37,19)
        56'b00000000000000000000000000001000001100000100010001110110,
        //Tile 798 (38,19)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 799 (39,19)
        56'b00000000000000000000000000001000000100001100010001101100,
        //Tile 800 (0,20)
        56'b00000000000000000000000000000000000000101000001001110111,
        //Tile 801 (1,20)
        56'b00000000000000000000000000000000000000001000101001111000,
        //Tile 802 (2,20)
        56'b00000000000000000000000000000000101000010000001001111001,
        //Tile 803 (3,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 804 (4,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 805 (5,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 806 (6,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 807 (7,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 808 (8,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 809 (9,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 810 (10,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 811 (11,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 812 (12,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 813 (13,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 814 (14,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 815 (15,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 816 (16,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 817 (17,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 818 (18,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 819 (19,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 820 (20,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 821 (21,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 822 (22,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 823 (23,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 824 (24,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 825 (25,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 826 (26,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 827 (27,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 828 (28,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 829 (29,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 830 (30,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 831 (31,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 832 (32,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 833 (33,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 834 (34,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 835 (35,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 836 (36,20)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 837 (37,20)
        56'b00000000000000000000000000000000000000101000001001110111,
        //Tile 838 (38,20)
        56'b00000000000000000000000000000000000000001000101001111000,
        //Tile 839 (39,20)
        56'b00000000000000000000000000000000101000010000001001111001,
        //Tile 840 (0,21)
        56'b00000000000000000000000000000001000000101000001001111011,
        //Tile 841 (1,21)
        56'b00000000000000000000000000000000000000001000101001111000,
        //Tile 842 (2,21)
        56'b00000000000000000000000000000001000000101000001001111100,
        //Tile 843 (3,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 844 (4,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 845 (5,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 846 (6,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 847 (7,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 848 (8,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 849 (9,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 850 (10,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 851 (11,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 852 (12,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 853 (13,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 854 (14,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 855 (15,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 856 (16,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 857 (17,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 858 (18,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 859 (19,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 860 (20,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 861 (21,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 862 (22,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 863 (23,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 864 (24,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 865 (25,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 866 (26,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 867 (27,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 868 (28,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 869 (29,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 870 (30,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 871 (31,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 872 (32,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 873 (33,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 874 (34,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 875 (35,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 876 (36,21)
        56'b00000000000000000000000000000001000000101000001001111101,
        //Tile 877 (37,21)
        56'b00000000000000000000000000000001000000101000001001111011,
        //Tile 878 (38,21)
        56'b00000000000000000000000000000000000000001000101001111000,
        //Tile 879 (39,21)
        56'b00000000000000000000000000000001000000101000001001111100,
        //Tile 880 (0,22)
        56'b00000000000000000000000000000001000000101000001001111110,
        //Tile 881 (1,22)
        56'b00000000000000000000000000000000000000001000101001111000,
        //Tile 882 (2,22)
        56'b00000000000000000000000000000001000000101000001001111111,
        //Tile 883 (3,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 884 (4,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 885 (5,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 886 (6,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 887 (7,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 888 (8,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 889 (9,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 890 (10,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 891 (11,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 892 (12,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 893 (13,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 894 (14,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 895 (15,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 896 (16,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 897 (17,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 898 (18,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 899 (19,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 900 (20,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 901 (21,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 902 (22,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 903 (23,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 904 (24,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 905 (25,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 906 (26,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 907 (27,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 908 (28,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 909 (29,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 910 (30,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 911 (31,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 912 (32,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 913 (33,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 914 (34,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 915 (35,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 916 (36,22)
        56'b00000000000000000000000000000000101001000000001010000000,
        //Tile 917 (37,22)
        56'b00000000000000000000000000000001000000101000001001111110,
        //Tile 918 (38,22)
        56'b00000000000000000000000000000000000000001000101001111000,
        //Tile 919 (39,22)
        56'b00000000000000000000000000000001000000101000001001111111,
        //Tile 920 (0,23)
        56'b00000000000000000000000000000000000000101000001010000001,
        //Tile 921 (1,23)
        56'b00000000000000000000000000000000000000101000001010000010,
        //Tile 922 (2,23)
        56'b00000000000000000000000000000000000000101000001010000011,
        //Tile 923 (3,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 924 (4,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 925 (5,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 926 (6,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 927 (7,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 928 (8,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 929 (9,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 930 (10,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 931 (11,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 932 (12,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 933 (13,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 934 (14,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 935 (15,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 936 (16,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 937 (17,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 938 (18,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 939 (19,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 940 (20,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 941 (21,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 942 (22,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 943 (23,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 944 (24,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 945 (25,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 946 (26,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 947 (27,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 948 (28,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 949 (29,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 950 (30,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 951 (31,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 952 (32,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 953 (33,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 954 (34,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 955 (35,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 956 (36,23)
        56'b00000000000000000000000000000000000000101000001001111010,
        //Tile 957 (37,23)
        56'b00000000000000000000000000000000000000101000001010000001,
        //Tile 958 (38,23)
        56'b00000000000000000000000000000000000000101000001010000010,
        //Tile 959 (39,23)
        56'b00000000000000000000000000000000000000101000001010000011,
        //Tile 960 (0,24)
        56'b00000000000000000000000000001100000100010000001010000100,
        //Tile 961 (1,24)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 962 (2,24)
        56'b00000000000000000000000000001100000100001000010010000101,
        //Tile 963 (3,24)
        56'b00000000000000000000000000000000000000101000001010000110,
        //Tile 964 (4,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 965 (5,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 966 (6,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 967 (7,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 968 (8,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 969 (9,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 970 (10,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 971 (11,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 972 (12,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 973 (13,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 974 (14,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 975 (15,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 976 (16,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 977 (17,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 978 (18,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 979 (19,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 980 (20,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 981 (21,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 982 (22,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 983 (23,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 984 (24,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 985 (25,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 986 (26,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 987 (27,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 988 (28,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 989 (29,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 990 (30,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 991 (31,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 992 (32,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 993 (33,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 994 (34,24)
        56'b00000000000000000000000000000000000000101000001010000111,
        //Tile 995 (35,24)
        56'b00000000000000000000000000000000000000101000001010001000,
        //Tile 996 (36,24)
        56'b00000000000000000000000000000000000000101000001010001001,
        //Tile 997 (37,24)
        56'b00000000000000000000000000001100000100010000001010000100,
        //Tile 998 (38,24)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 999 (39,24)
        56'b00000000000000000000000000001100000100001000010010000101,
        //Tile 1000 (0,25)
        56'b00000000000000000000000000001000001100000100010010001010,
        //Tile 1001 (1,25)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1002 (2,25)
        56'b00000000000000000000000000001000001100000100010010010011,
        //Tile 1003 (3,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1004 (4,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1005 (5,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1006 (6,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1007 (7,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1008 (8,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1009 (9,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1010 (10,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1011 (11,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1012 (12,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1013 (13,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1014 (14,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1015 (15,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1016 (16,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1017 (17,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1018 (18,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1019 (19,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1020 (20,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1021 (21,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1022 (22,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1023 (23,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1024 (24,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1025 (25,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1026 (26,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1027 (27,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1028 (28,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1029 (29,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1030 (30,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1031 (31,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1032 (32,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1033 (33,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1034 (34,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1035 (35,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1036 (36,25)
        56'b00000000000000000000000000001000001100000100010000111000,
        //Tile 1037 (37,25)
        56'b00000000000000000000000000001100000100010000001010001110,
        //Tile 1038 (38,25)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1039 (39,25)
        56'b00000000000000000000000000001100000100010000001010001110,
        //Tile 1040 (0,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1041 (1,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1042 (2,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1043 (3,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1044 (4,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1045 (5,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1046 (6,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1047 (7,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1048 (8,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1049 (9,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1050 (10,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1051 (11,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1052 (12,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1053 (13,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1054 (14,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1055 (15,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1056 (16,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1057 (17,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1058 (18,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1059 (19,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1060 (20,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1061 (21,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1062 (22,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1063 (23,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1064 (24,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1065 (25,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1066 (26,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1067 (27,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1068 (28,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1069 (29,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1070 (30,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1071 (31,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1072 (32,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1073 (33,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1074 (34,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1075 (35,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1076 (36,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1077 (37,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1078 (38,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1079 (39,26)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1080 (0,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1081 (1,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1082 (2,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1083 (3,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1084 (4,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1085 (5,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1086 (6,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1087 (7,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1088 (8,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1089 (9,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1090 (10,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1091 (11,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1092 (12,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1093 (13,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1094 (14,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1095 (15,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1096 (16,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1097 (17,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1098 (18,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1099 (19,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1100 (20,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1101 (21,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1102 (22,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1103 (23,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1104 (24,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1105 (25,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1106 (26,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1107 (27,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1108 (28,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1109 (29,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1110 (30,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1111 (31,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1112 (32,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1113 (33,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1114 (34,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1115 (35,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1116 (36,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1117 (37,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1118 (38,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1119 (39,27)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1120 (0,28)
        56'b00000000000000000000100100100000011000010100011110010100,
        //Tile 1121 (1,28)
        56'b00000000000000000000000000100100011000100000010110010101,
        //Tile 1122 (2,28)
        56'b00000000000000000000000000100100011000100000010110010101,
        //Tile 1123 (3,28)
        56'b00000000000000000000100100011000100000011100010110010110,
        //Tile 1124 (4,28)
        56'b00000000000000000000000001011101011001010101010010010111,
        //Tile 1125 (5,28)
        56'b00000000000000000000000001011101011001010101010010011000,
        //Tile 1126 (6,28)
        56'b00000000000000000000000001011101011001010101010010011000,
        //Tile 1127 (7,28)
        56'b00000000000000000000000001011101011001010101010010011000,
        //Tile 1128 (8,28)
        56'b00000000000000000000000001011101011001010101010010011001,
        //Tile 1129 (9,28)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1130 (10,28)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1131 (11,28)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1132 (12,28)
        56'b10100110100010011100010010011000001100001000000110011010,
        //Tile 1133 (13,28)
        56'b00000000000010011010011100010000001100001000000110011011,
        //Tile 1134 (14,28)
        56'b00000000000010011100010010011000001100001000000110011100,
        //Tile 1135 (15,28)
        56'b00000000000000010010011110011000001100001000000110011101,
        //Tile 1136 (16,28)
        56'b00000000000000000000010010011000001100001000000110011110,
        //Tile 1137 (17,28)
        56'b00000000000000000000010010011000001100001000000110011111,
        //Tile 1138 (18,28)
        56'b00000000000010011100010010011000001100001000000110100000,
        //Tile 1139 (19,28)
        56'b00000000000000000010011110011000001100001000000110100001,
        //Tile 1140 (20,28)
        56'b00000010100010100110011000010000001100001000000110100010,
        //Tile 1141 (21,28)
        56'b00000000000000000000010010011000001100001000000110100011,
        //Tile 1142 (22,28)
        56'b00000000000000000010011000010000001100001000000110100100,
        //Tile 1143 (23,28)
        56'b00000000000000000000000010011000001100001000000110100101,
        //Tile 1144 (24,28)
        56'b00000000000000000000000010011000001100001000000110100110,
        //Tile 1145 (25,28)
        56'b00000000000000000010100000010000001100001000000110100111,
        //Tile 1146 (26,28)
        56'b00000000000000000010100000010000001100001000000110101000,
        //Tile 1147 (27,28)
        56'b00000000000000000000100100100000011000010100011110010100,
        //Tile 1148 (28,28)
        56'b00000000000000000000000000100100011000100000010110010101,
        //Tile 1149 (29,28)
        56'b00000000000000000000000000100100011000100000010110010101,
        //Tile 1150 (30,28)
        56'b00000000000000000000000000100100011000100000010110010101,
        //Tile 1151 (31,28)
        56'b00000000000000000000100100011000100000011100010110010110,
        //Tile 1152 (32,28)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1153 (33,28)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1154 (34,28)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1155 (35,28)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1156 (36,28)
        56'b00000000000000000000000000000000001100001000000100001000,
        //Tile 1157 (37,28)
        56'b00000000000000000000000100101000001100010000001010101001,
        //Tile 1158 (38,28)
        56'b00000000000000000000000100001100101000001000010010101010,
        //Tile 1159 (39,28)
        56'b00000000000000000000000100001100101000001000010010101011,
        //Tile 1160 (0,29)
        56'b00000000000000000000000000000000000000011000010110101100,
        //Tile 1161 (1,29)
        56'b00000000000000000000000000001100000100010000001010101101,
        //Tile 1162 (2,29)
        56'b00000000000000000000000000000000000000000000011010101110,
        //Tile 1163 (3,29)
        56'b00000000000000000000000000000000000000010100011010101111,
        //Tile 1164 (4,29)
        56'b00000000000000000000000001010001011101011001010110110000,
        //Tile 1165 (5,29)
        56'b00000000000000000000000001010101011101011001010010110001,
        //Tile 1166 (6,29)
        56'b00000000000000000000000001010101011101011001010010110001,
        //Tile 1167 (7,29)
        56'b00000000000000000000000001010101011101011001010010110001,
        //Tile 1168 (8,29)
        56'b00000000000000000000000001010101011101011001010010110010,
        //Tile 1169 (9,29)
        56'b00000000000000000000000000001100000100010000001010110011,
        //Tile 1170 (10,29)
        56'b00000000000000000000000000001100001000000100010010110100,
        //Tile 1171 (11,29)
        56'b00000000000000000000000000001100000100001000010010110101,
        //Tile 1172 (12,29)
        56'b00000000000000001110011110101010100010100100010010110110,
        //Tile 1173 (13,29)
        56'b00000000000010100100010010101010100010011010011110110111,
        //Tile 1174 (14,29)
        56'b00000000000000000010100110100000010010011010011110111000,
        //Tile 1175 (15,29)
        56'b00000000000000000010100110100000010010011110011010111001,
        //Tile 1176 (16,29)
        56'b00000010100010100110011010011100001000000100010010111010,
        //Tile 1177 (17,29)
        56'b00000010100110100010011010011100010000001000000110111011,
        //Tile 1178 (18,29)
        56'b00000000000000000010100110100010011110011000010010111100,
        //Tile 1179 (19,29)
        56'b00000000000000000010100010100100010010011110011010111101,
        //Tile 1180 (20,29)
        56'b00000000000000000010011110100000010010100110011010111110,
        //Tile 1181 (21,29)
        56'b00000000000000000010100010011110100110011000010010111111,
        //Tile 1182 (22,29)
        56'b00000000000000000010011110100010100110011000010011000000,
        //Tile 1183 (23,29)
        56'b00000000000000000010100110100010011100010010011011000001,
        //Tile 1184 (24,29)
        56'b00000000010010011100000100001010100010100110011011000010,
        //Tile 1185 (25,29)
        56'b00000000000010011010011110100110100000010000000111000011,
        //Tile 1186 (26,29)
        56'b00000000000000000000000000000000000000010010100111000100,
        //Tile 1187 (27,29)
        56'b00000000000000000000000000000000000000011000010110101100,
        //Tile 1188 (28,29)
        56'b00000000000000000000000000000000000000000000011010101110,
        //Tile 1189 (29,29)
        56'b00000000000000000000000000000000000000000000011010101110,
        //Tile 1190 (30,29)
        56'b00000000000000000000000000000000000000000000011010101110,
        //Tile 1191 (31,29)
        56'b00000000000000000000000000000000000000010100011010101111,
        //Tile 1192 (32,29)
        56'b00000000000000000000000001101101101001100101100011000101,
        //Tile 1193 (33,29)
        56'b00000000000000000000000000000001101101101001100111000110,
        //Tile 1194 (34,29)
        56'b00000000000000000000000000000001101101101001100111000110,
        //Tile 1195 (35,29)
        56'b00000000000000000000000000000001101101101001100111000110,
        //Tile 1196 (36,29)
        56'b00000000000000000000000001101101101001100001100111000111,
        //Tile 1197 (37,29)
        56'b00000000000000000000000000101000001100000100010011001000,
        //Tile 1198 (38,29)
        56'b00000000000000000000000000000000001100000100101011001001,
        //Tile 1199 (39,29)
        56'b00000000000000000000000000010000001100000100101011001010
    };

    assign data = ROM[addr];

endmodule