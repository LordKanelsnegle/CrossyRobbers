module tile_rom (
    input logic [11:0] addr,
    output logic [47:0] data
);

    parameter bit [47:0] ROM [3248] = '{
        //tile_code 0
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011011011011011011011011011011011011011011011,
        //tile_code 1
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b001001001001001001001001001001001001001011000010,
        48'b000000000000000000000000000000000000000000000010,
        48'b001001001001001001001001001001001001001001001010,
        48'b011011011011011011011011011011011011011011011010,
        48'b010010010010010010010010010010010010010010010001,
        //tile_code 2
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001010000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000011011011011011011011011011011011011011011011,
        48'b000000000000000000000000000000000000000000000000,
        48'b000100100100100100100100100100100100100100100100,
        48'b000100100100100100100100100100100100100100100100,
        48'b000100100100100100100100100100100100100100100100,
        48'b000100100100100100100100100100100100100100100100,
        48'b000100100100100100100100100100100100100100100100,
        48'b000100100100100100100100100100100100100100100100,
        48'b010000000000000000000000000000000000000000000000,
        //tile_code 3
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b001001001001001001001001001001001001001001001001,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b001001001001001001001001001001001001001001001001,
        //tile_code 4
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b001001001001001001001001001001001001010000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b011011011011011011011011011011011011011011011001,
        48'b001001001001001001001001001001001001001001001001,
        48'b100100100100100100100100100100100100100100100001,
        48'b100100100100100100100100100100100100100100100001,
        48'b100100100100100100100100100100100100100100100001,
        48'b100100100100100100100100100100100100100100100001,
        48'b100100100100100100100100100100100100100100100001,
        48'b100100100100100100100100100100100100100100100001,
        48'b001001001001001001001001001001001001001001001010,
        //tile_code 5
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000010010010011010010010011010010010011010010010,
        48'b000010010010010010010010010010010010010010010010,
        48'b100100100000000100100000000100100000000100100000,
        //tile_code 6
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000010010010000010010010000010010010000010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b011100100011011100100011011100100011011100100011,
        //tile_code 7
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000010010010000010010010000010010010000010010011,
        48'b010010010010010010010010010010010010010010010011,
        48'b011100100011011100100011011100100011011100100100,
        //tile_code 8
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        //tile_code 9
        48'b000000001010011010011010011010011010011001100001,
        48'b000000001010011010011010011010011010011001100001,
        48'b000000001010011010011010011010011010011001100001,
        48'b101101001010011010011010011010011010011001100001,
        48'b000000001010011010011010011010011010011001100001,
        48'b000000001010011010011010011010011010011001100001,
        48'b000000001010011010011010011010011010011110001110,
        48'b101101001010011010011010011010011010011001000001,
        48'b000000001001001001001001001001001001001001001001,
        48'b000000001000000000000000000000000000000001110001,
        48'b000000110001001001001001001001001001001110110001,
        48'b101101001110110110110110110110110110110110110001,
        48'b000000001110001001001001001001001001001001110001,
        48'b000000001001110001001001001001001001001110001001,
        48'b000000001001110110001001001001001001110110001001,
        48'b101101001001001001001001001001001001001001001001,
        //tile_code 10
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000010010010010010010010010010010010010010010000,
        48'b000010011011011011011011011011011011011011010000,
        //tile_code 11
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000001010010001000000000,
        48'b000000011000000000000000001010100100010001001000,
        48'b000000000000000000001001001010100100010001011001,
        48'b011000000000000001011011001010001001010001000001,
        48'b000000000000000001000000000001000001001001001000,
        48'b000000000000000000001001001001001000000000000000,
        48'b000000000000101101000000000011000000000000000000,
        48'b000000000101110110101000000000000000000000000000,
        48'b011000101110100100110101000000000000000000000000,
        48'b000101110110100100110110101000000000000000000000,
        48'b000101110101110110101110101001001000000000000000,
        48'b000001101101110110101101011011011001000000000000,
        48'b001011011000101101001001000000001000000011000000,
        48'b001000000000001000000000001001000011011011000000,
        48'b000001001001000000000000000000000011011000000000,
        //tile_code 12
        48'b000001001001001001001010010010010010010010010010,
        48'b000001001001001001001001010010010010010010010010,
        48'b000001001001001001001001001010010010010010010011,
        48'b001000001001001001001001001010010010010010010011,
        48'b010001000011001001001011001001010010010010010010,
        48'b001001000001011011011001011001001010010010010010,
        48'b001001000001001001001001001011001010010010010010,
        48'b001001000001001001001001001001011001010010010010,
        48'b001001000001001001001001001001001011011011011010,
        48'b010001000001011001001001001001001001001001001011,
        48'b001001001000011001001001001001001001001001001001,
        48'b001001001001011011011011011001001001001001001001,
        48'b001001001001001000000011011011001001001001001001,
        48'b001001001001001010001000011011011011001001011001,
        48'b001001001001001001001001000011011011011011011001,
        48'b001001001001001001001001001000011011011011011011,
        //tile_code 13
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b010010010010001000000000000000000000000000000001,
        48'b000000000000010010010000000000000000000001010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000001000000000001,
        48'b000010010000000001000000000000001001001001001001,
        48'b010001001010010001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001010010010010,
        48'b010001001001001001001001001001001010001001001001,
        //tile_code 14
        48'b000000000000000000000001010010001010010010011010,
        48'b000000000000000000001010001001010010010010010011,
        48'b000000000000000010001010010010010010010010010011,
        48'b000000001000001001010010010010010010010010001011,
        48'b010001010001010010010010010010010010010001001011,
        48'b001010010010010010010010010010010010001001001011,
        48'b000010010010010010010010010010001001001001001011,
        48'b010010010010010010010010010001001001001001001011,
        48'b010010010010010010001010001001001001001001011010,
        48'b010010010010010010001001001001001001001011010010,
        48'b010010010010010010001001001001001001011010010010,
        48'b010010010010010001001001001011011011010010010010,
        48'b010001010010001001001001011010010010010010010010,
        48'b001010010001001001001011010010010010010000010010,
        48'b010010001001001001011010010010010000000000010010,
        48'b010001001001001011010010010010010000000010010010,
        //tile_code 15
        48'b000001000010011010011010011010011010011000100100,
        48'b000001000010011010011010011010011010011000100100,
        48'b000001000010011010011010011010011010011000100100,
        48'b000001000010011010011010011010011010011000101101,
        48'b000001000010011010011010011010011010011000100110,
        48'b000001000010011010011010011010011010011000100110,
        48'b110000110010011010011010011010011010011000100110,
        48'b000100000010011010011010011010011010011000101101,
        48'b000000000000000000000000000000000000000000100100,
        48'b000110000100100100100100100100100100100000100100,
        48'b000110110000000000000000000000000000000110100100,
        48'b000110110110110110110110110110110110110000101101,
        48'b000110000000000000000000000000000000110000100110,
        48'b000000110000000000000000000000000110000000100110,
        48'b000000110110000000000000000000110110000000100110,
        48'b000000000000000000000000000000000000000000101101,
        //tile_code 16
        48'b000001001000000001001000000001001000000001001000,
        48'b001010011001001010011001001010011001001010011001,
        48'b001001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b001010011000000010011000000010011000000010011000,
        48'b001010011000000010011000000010011000000010011000,
        48'b001001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b001010011000000010011000000010011000000010011000,
        48'b001010011000000010011000000010011000000010011000,
        48'b001001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b001010011000000010011000000010011000000010011000,
        48'b001010011000000010011000000010011000000010011000,
        48'b001001001000000001001000000001001000000001001000,
        48'b001001001001001001001001001001001001001001001001,
        //tile_code 17
        48'b000001001000000001001000000001001000000001001000,
        48'b001010011001001010011001001010011001001010011001,
        48'b000001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011000,
        48'b000010011000000010011000000010011000000010011000,
        48'b000001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011000,
        48'b000010011000000010011000000010011000000010011000,
        48'b000001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011000,
        48'b000010011000000010011000000010011000000010011000,
        48'b000001001000000001001000000001001000000001001000,
        48'b001001001001001001001001001001001001001001001001,
        //tile_code 18
        48'b000001001000000001001000000001001000000001001000,
        48'b001010011001001010011001001010011001001010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001001001001001001001001001001001001001001001001,
        //tile_code 19
        48'b000001001001001001001001001001001001001001001001,
        48'b001010010010010010010010010010010010010010010010,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001000001000001000001000001000001000001000001000,
        48'b000001001001001001001001001001001001001001001001,
        //tile_code 20
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000011000011000011000011000011000011000011000011,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 21
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001000001000001000001000001000001000001000000,
        48'b000000000000000000000000000000000000000000000001,
        //tile_code 22
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        //tile_code 23
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        //tile_code 24
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010001010010010010010010010010010010010010,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010010010010010010010010010001010010010010,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010010010001010010010010010010010010010010,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010010010010010010010010001010010010010010,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 25
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001000001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001000001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001000001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001000001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        //tile_code 26
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010000010010010010010010010010010010010001,
        48'b000000000000000000000000000000000000000000000001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010000010010010001,
        48'b000000000000000000000000000000000000000000000001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010000010010010010010010010010010001,
        48'b000000000000000000000000000000000000000000000001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010000010010010010001,
        48'b000000000000000000000000000000000000000000000001,
        48'b001001001001001001001001001001001001001001001001,
        //tile_code 27
        48'b000001001000001001001001001001001000001001001001,
        48'b000010010000010010010010010010010000010010010010,
        48'b000010010000010010010010010010010000010010010010,
        48'b000011011011011011011011011011011011011011011011,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011011,
        48'b000001001000001001001001001001001000001001001001,
        48'b000010010000010010010010010010010000010010010010,
        48'b000010010000010010010010010010010000010010010010,
        48'b000011011011011011011011011011011011011011011011,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011011,
        //tile_code 28
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010001010010010010010010010001010010010010,
        48'b010010010001010010010010010010010001010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010001010010010010010010010001010010010010,
        48'b010010010001010010010010010010010001010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011011,
        //tile_code 29
        48'b000000000001000000000000000000000001000000000001,
        48'b010010010001010010010010010010010001010010010001,
        48'b010010010001010010010010010010010001010010010001,
        48'b011011011011011011011011011011011011011011011001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011001,
        48'b000000000001000000000000000000000001000000000001,
        48'b010010010001010010010010010010010001010010010001,
        48'b010010010001010010010010010010010001010010010001,
        48'b011011011011011011011011011011011011011011011001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011001,
        //tile_code 30
        48'b000000000001000000000000000000000001000001010001,
        48'b000000000001000000000000000000000001000010000010,
        48'b000000000001000000000000000000000001000010010010,
        48'b011011011011011011011011011011011011011010100010,
        48'b000000001010010010010010010010010010010010100010,
        48'b000000010000000000000000000000000000000010100010,
        48'b000000010010010010010010010010010010010010100010,
        48'b011011010101110101110101110101110101110010100010,
        48'b000000010101110101110101110101110101110010100010,
        48'b000000010101110101110101110101110101110010100010,
        48'b000000010101110101110101110101110101110010100010,
        48'b011011010101110101110101110101110101110010100010,
        48'b000000010101110101110101110101110101110010100010,
        48'b000000010101110101110101110101110101110010100010,
        48'b000000010101110101110101110101110101110010100010,
        48'b011011010101110101110101110101110101110010100010,
        //tile_code 31
        48'b000000000000000000000000000000001001010010010010,
        48'b000000000000000000000000000000000000001001001001,
        48'b000000011000000000000000000000000000000000011000,
        48'b000000000000000000000000000000000000000000011011,
        48'b011000000000000011000000000000000000000000000011,
        48'b000000000000000011011011000000000000000000000000,
        48'b000000000000000000011011000000011000000000000000,
        48'b000000000000100100000000000011000000000000000000,
        48'b000000000100101101100000000000000000000000000000,
        48'b011000100101110110101100000000000000000000000000,
        48'b000100101101110110101101100000000000000000000000,
        48'b000100101100101101100101100001001000000000000000,
        48'b000001100100101101100100011011011001000000000000,
        48'b001011011000100100001001000000001000000011000000,
        48'b001000000000001000000000001001000011011011000000,
        48'b000001001001000000000000000000000011011000000000,
        //tile_code 32
        48'b000000000001001001001000000000000001001001001001,
        48'b010000000000000000001001001000001001001001000000,
        48'b010000000000000000000000000000000000000000000000,
        48'b001010000000010010000000000000000000000000010010,
        48'b011001010010100101010010000000000000000010001011,
        48'b001001001001100101101101010010010010010001001001,
        48'b001001001001100101101101101101101100001001001001,
        48'b001001001001100101101101101101101100001001001001,
        48'b001001001001100110101101101101110100001001001001,
        48'b011001100100110110110110110110110110100001001001,
        48'b100100101101110100100110100100110110110100001001,
        48'b100100100100100001100110100100100100101101100001,
        48'b001001001001001001100110100001001001100100001001,
        48'b001001001001001011100101100001001001001011001001,
        48'b001001001001001001100101100001001011011011001001,
        48'b001001001001001001001100001001001011011001001001,
        //tile_code 33
        48'b000000001001001010010010010010001001010010010010,
        48'b000001010010010010010010010001011011001010010010,
        48'b001010100010010010010010001011101101011001001010,
        48'b010010010010010010001001001011101101011001100001,
        48'b100010010010010001100100001011001001011001010001,
        48'b010010010010010001010010010001010001001001001010,
        48'b010010010010010010001001001001001010010010010010,
        48'b010010010010010010010010010100010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b100010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010100010010010010010010010100010010,
        48'b010010010010010010010010010010010100100100010010,
        48'b010010010010010010010010010010010100100010010010,
        //tile_code 34
        48'b000001000000010010010010010010010000010010010010,
        48'b001010001000010010010010010010010000010010010010,
        48'b001001001000010010010010010010010000010010010010,
        48'b001011001100100100100100100100100100100100100100,
        48'b001011001001001001001001001001001001001000010000,
        48'b001011001010010010010010010010010010010001010000,
        48'b001011001001001001001001001001001001001001010000,
        48'b001011001101110101110101110101110101110001100100,
        48'b001011001101110101110101110101110101110001010010,
        48'b001011001101110101110101110101110101110001010010,
        48'b001011001101110101110101110101110101110001010010,
        48'b001011001101110101110101110101110101110001100100,
        48'b001011001101110101110101110101110101110001010000,
        48'b001011001101110101110101110101110101110001010000,
        48'b001011001101110101110101110101110101110001010000,
        48'b001011001101110101110101110101110101110001100100,
        //tile_code 35
        48'b000001001000001001001001001001001000001001001001,
        48'b000010010000010010010010010010010000010010010010,
        48'b000010010000010010010010010010010000010010010010,
        48'b000011011011011011011011011011011011011011011011,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011011,
        48'b000001001000001001001001001001001000001001001001,
        48'b000010010000010010010010010010010000010010010010,
        48'b000010010000010010010010010010010000010010010010,
        48'b000011011011011011011011011011011011011011011011,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011011,
        //tile_code 36
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010001010010010010010010010001010010010010,
        48'b010010010001010010010010010010010001010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010001010010010010010010010001010010010010,
        48'b010010010001010010010010010010010001010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011011,
        //tile_code 37
        48'b000000000001000000000000000000000001000000000001,
        48'b010010010001010010010010010010010001010010010001,
        48'b010010010001010010010010010010010001010010010001,
        48'b011011011011011011011011011011011011011011011001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011001,
        48'b000000000001000000000000000000000001000000000001,
        48'b010010010001010010010010010010010001010010010001,
        48'b010010010001010010010010010010010001010010010001,
        48'b011011011011011011011011011011011011011011011001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011001,
        //tile_code 38
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001011011011011011011011011011011011001001,
        48'b000100100011011011011011011011011011001011100100,
        48'b000100100011011011011011011011011001001011100100,
        48'b000100100011011011011011011011001001011011100100,
        48'b000100100011011011011011011001001011011011100100,
        48'b000100100011011011011011001001011011011011100100,
        48'b000100100011011011011001001011011011011011100100,
        48'b000100100011011011001001011011011011001011100100,
        48'b000100100011011001001011011011011001011011100100,
        48'b000100100011001001011011011011001011011011100100,
        48'b000100100011001011011011011001011011011011100100,
        //tile_code 39
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001011011011011011011011011011011011001001,
        48'b100100100011011011011011011011011011001011100100,
        48'b100100100011011011011011011011011001001011100100,
        48'b100100100011011011011011011011001001011011100100,
        48'b100100100011011011011011011001001011011011100100,
        48'b100100100011011011011011001001011011011011100100,
        48'b100100100011011011011001001011011011011011100100,
        48'b100100100011011011001001011011011011001011100100,
        48'b100100100011011001001011011011011001011011100100,
        48'b100100100011001001011011011011001011011011100100,
        48'b100100100011001011011011011001011011011011100100,
        //tile_code 40
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 41
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 42
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001011011011011011011011011011011011001000,
        48'b100100100011011011011011011011011011001011100000,
        48'b100100100011011011011011011011011001001011100000,
        48'b100100100011011011011011011011001001011011100000,
        48'b100100100011011011011011011001001011011011100000,
        48'b100100100011011011011011001001011011011011100000,
        48'b100100100011011011011001001011011011011011100000,
        48'b100100100011011011001001011011011011001011100000,
        48'b100100100011011001001011011011011001011011100000,
        48'b100100100011001001011011011011001011011011100000,
        48'b100100100011001011011011011001011011011011100000,
        //tile_code 43
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001010010001001010010001001010010001001000,
        48'b000001001010010001001010010001001010010001001000,
        48'b000001001010010001001010010001001010010001001000,
        48'b000011011100100011011100100011011100100011011000,
        48'b000000000101101000000101101000000101101000000000,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101011101000000000000011011000000000011101011101,
        48'b101011101000000000011011000000000011000101011101,
        48'b101011101000000011011000000000011000000101011101,
        48'b101011101000011011000000000011000000000101011101,
        48'b101011000101101101101101101101101101101000011101,
        48'b101011000110110110110110110110110110110000011101,
        48'b101011011011011011011011011011011011011011011101,
        48'b000101101101101101101101101101101101101101101000,
        //tile_code 44
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001011011011011011011011011011011011001001000,
        48'b100100011011011011011011011011011001011100100000,
        48'b100100011011011011011011011011001001011100100000,
        48'b100100011011011011011011011001001011011100100000,
        48'b100100011011011011011011001001011011011100100000,
        48'b100100011011011011011001001011011011011100100000,
        48'b100100011011011011001001011011011011011100100000,
        48'b100100011011011001001011011011011001011100100000,
        48'b100100011011001001011011011011001011011100100000,
        48'b100100011001001011011011011001011011011100100000,
        48'b100100011011011011011011011011011011011100100000,
        //tile_code 45
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000001001001001001001001010010001001001000000,
        48'b000000001001001001001001010010001001001001000000,
        48'b000000011011011011011010010011011011011011000000,
        48'b000000011011011011010010011011011011011011000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000001001001001001001001010001001001001000000,
        48'b000000001001001001001001010001001001001001000000,
        48'b000000001001001001001010001001001001001001000000,
        48'b000000001001001001010001001001001001001001000000,
        48'b000000001001001010001001001001001001001001000000,
        48'b000000001001010001001001001001001001001001000000,
        48'b000000001010001001001001001001001001001001000000,
        48'b000000010001001001001001001011001001001011000000,
        //tile_code 46
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000001001001001001001001010010001001001000000,
        48'b000000001001001001001001010010001001001001000000,
        48'b000000011011011011011010010011011011011011000000,
        48'b000000011011011011010010011011011011011011000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000001001001001001001001010001001001001000000,
        48'b000000001001001001001001010001001001001001000000,
        48'b000000001001001001001010001001001001001001000000,
        48'b000000001001001001010001001001001001001001000000,
        48'b000000001001001010001001001001001001001001000000,
        48'b000000001001010001001001001001001001001001000000,
        48'b000000001010001001001001001001001001001001000000,
        48'b000000011001001001011001001001001001001001000000,
        //tile_code 47
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001011011011011011011011011011011011001001,
        48'b000100100011011011011011011011011011001011100100,
        48'b000100100011011011011011011011011001001011100100,
        48'b000100100011011011011011011011001001011011100100,
        48'b000100100011011011011011011001001011011011100100,
        48'b000100100011011011011011001001011011011011100100,
        48'b000100100011011011011001001011011011011011100100,
        48'b000100100011011011001001011011011011001011100100,
        48'b000100100011011001001011011011011001011011100100,
        48'b000100100011001001011011011011001011011011100100,
        48'b000100100011011011011011011011011011011011100100,
        //tile_code 48
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001011011011011011011011011011011011001000,
        48'b100100100011011011011011011011011011001011100000,
        48'b100100100011011011011011011011011001001011100000,
        48'b100100100011011011011011011011001001011011100000,
        48'b100100100011011011011011011001001011011011100000,
        48'b100100100011011011011011001001011011011011100000,
        48'b100100100011011011011001001011011011011011100000,
        48'b100100100011011011001001011011011011001011100000,
        48'b100100100011011001001011011011011001011011100000,
        48'b100100100011001001011011011011001011011011100000,
        48'b100100100011011011011011011011011011011011100000,
        //tile_code 49
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001010010001001010010001001010010001001010,
        48'b000001001010010001001010010001001010010001001010,
        48'b000001001010010001001010010001001010010001001010,
        48'b000011011100100011011100100011011100100011011100,
        48'b000000000101101000000101101000000101101000000101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101011101000011000000000000000000011000101011101,
        48'b101011101011000000000000000000011000000101011101,
        48'b101011101000000000000000000011000000000101011101,
        48'b101011101000000000000000011000000000000101011101,
        48'b101011101000000000000011000000000000000101011101,
        48'b101011101000000000011000000000000000000101011101,
        48'b101000101101101101101101101101101101101101000101,
        48'b101101011011011011011011011011011011011011101101,
        //tile_code 50
        48'b000000000000000000000000000000000000000000000000,
        48'b001010010001001010010001001010010001001010010000,
        48'b001010010001001010010001001010010001001010010000,
        48'b001010010001001010010001001010010001001010010000,
        48'b011100100011011100100011011100100011011100100000,
        48'b101000000101101000000101101000000101101000000000,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101100101000100000000000000000000100000101100101,
        48'b101100101100000000000000000000100000000101100101,
        48'b101100101000000000000000000100000000000101100101,
        48'b101100101000000000000000100000000000000101100101,
        48'b101100101000000000000100000000000000000101100101,
        48'b101100101000000000100000000000000000000101100101,
        48'b101000101101101101101101101101101101101101000101,
        48'b101101100100100100100100100100100100100100101101,
        //tile_code 51
        48'b000000000000000000000000000000000000000000000000,
        48'b000001010010010010010010010010010010010010001000,
        48'b000001000000000000000000000000000000000000001000,
        48'b000001000011011011011011011011011011011000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000000000000000000000000000000000000001000,
        48'b000001000000000000000000000000000000000000001000,
        48'b000001001001001001001001001001001001100100001000,
        //tile_code 52
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010001011011011011011011011011011011011011001010,
        48'b010001001001001001001001001001001001001001001010,
        48'b010001100100100101100101100101100100100100001010,
        48'b010001100100100100101100101100101100100100001010,
        48'b010001100100110101110101110101100100100100001010,
        48'b010001100110010010010010010010110110100100001010,
        48'b010001100110110110110110110110111100110100001010,
        48'b010001100100111110110110110111100111100100001010,
        48'b010001100111111111111111111111111100100100001010,
        48'b010001100111110110110110110110111100100100001010,
        48'b010001100100111111111111111111100100100100001010,
        48'b010001001001001001001001001001001001001001001010,
        48'b000001000000000000000000000000000000000000001000,
        48'b001001001001001001001001001001001001001001001001,
        //tile_code 53
        48'b000001001000001001001001001001001000001001001000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000011011011011011011011011011011011011011011000,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011000,
        48'b000001001000001001001001001001001000001001001000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000011011011011011011011011011011011011011011000,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011000,
        //tile_code 54
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011011011011011011011011011011011011011011011,
        //tile_code 55
        48'b000001001001001001001001001001001001001001001010,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000010001001001001001001001001001001001001001011,
        48'b011000001001001001001001001001001001001001001011,
        48'b011000010001001001001001001001001001001001001011,
        48'b011011000010010001001001001001001001001001001011,
        48'b011011011000000010010010010010010010010010010010,
        48'b011011011011011000000000000000000000000000000000,
        //tile_code 56
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 57
        48'b000001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001000010,
        48'b001001001001001001001001001001001001001001010011,
        48'b001001001001001001001001001001001001001000010011,
        48'b001001001001001001001001001001001000000010011011,
        48'b000000000000000000000000000000000010010011011011,
        48'b010010010010010010010010010010010011011011011011,
        //tile_code 58
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010001011010011011011011011011011010011011001010,
        48'b010001001001001001001001001001001001001001001010,
        48'b010001100100100100100101100100100100100100001010,
        48'b010001100100100100100011101101100100100100001010,
        48'b010001100100100100100110011011101101100100001010,
        48'b010001100100100100110110110110011011101100001010,
        48'b010001100100100100110111111110110110011101001010,
        48'b010001100100100110110111111110111110011100001010,
        48'b010001100100110111110110110110101011100100001010,
        48'b010001100100110110110110101011100100100100001010,
        48'b010001100110110110101011100100100100100100001010,
        48'b010001001001001001001001001001001001001001001010,
        48'b000001000000000000000000000000000000000000001000,
        48'b001001001001001001001001001001001001001001001001,
        //tile_code 59
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001010010001001010010001001010010001001010,
        48'b000001001010010001001010010001001010010001001010,
        48'b000001001010010001001010010001001010010001001010,
        48'b000011000100100011000100100011000100100011000100,
        48'b000000011011011000011011011000011011011000011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b101110101111111111111111111101110110110110110101,
        48'b101110101111111111111111111101110101101101110101,
        48'b101110101111111111111111111101110101111101110101,
        48'b101110101111111111111111111101110101111101110101,
        48'b101110101111111111111111111101110101101101110101,
        48'b101110101111111111111111111101110111111111110101,
        48'b101110101111111111111111111101110101101101110101,
        48'b101110101111111111111111111101110101111101110101,
        //tile_code 60
        48'b000000000000000000000000000000000000000000000000,
        48'b001010010001001010010001001010010001001010010000,
        48'b001010010001001010010001001010010001001010010000,
        48'b001010010001001010010001001010010001001010010000,
        48'b011100000011011100000011011100000011011100000000,
        48'b100000100100100000100100100000100100100000100000,
        48'b100100100100100100100100100100100100100100100100,
        48'b100100100100100100100100100100100100100100100100,
        48'b101110110110110110101111111111111111111101110101,
        48'b101110101101101110101111111111111111111101110101,
        48'b101110101111101110101111111111111111111101110101,
        48'b101110101111101110101111111111111111111101110101,
        48'b101110101101101110101111111111111111111101110101,
        48'b101110111111111110101111111111111111111101110101,
        48'b101110101101101110101111111111111111111101110101,
        48'b101110101111101110101111111111111111111101110101,
        //tile_code 61
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001010010001001010010001001010010001001010,
        48'b000001001010010001001010010001001010010001001010,
        48'b000001001010010001001010010001001010010001001010,
        48'b000011011100100011011100100011011100100011011100,
        48'b000000000101101000000101101000000101101000000101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b110110000000000000011000000000000000000000000000,
        48'b110110000000000011000000000000000000000000000011,
        48'b110110000000011000000000000000000000000000011011,
        48'b110110000011000000000000000000000000000011011000,
        48'b110110011101101101101101101101101101011011101101,
        48'b110110101101101101101101101101101011011101101101,
        48'b110110110110110110110110110110110110110110110110,
        48'b110110110110110110110110110110110110110110110110,
        //tile_code 62
        48'b000000000000000000000000000000000000000000000000,
        48'b001010010001001010010001001010010001001010010000,
        48'b001010010001001010010001001010010001001010010000,
        48'b001010010001001010010001001010010001001010010000,
        48'b011100100011011100100011011100100011011100100000,
        48'b101000000101101000000101101000000101101000000000,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b100100000000000000000000100000000000000000110110,
        48'b100000000000000000000100000000000000000000110110,
        48'b000000000000000000100000000000000000000000110110,
        48'b000000000000000100000000000000000000000000110110,
        48'b101101101101100101101101101101101101101101110110,
        48'b101101101100101101101101101101101101101101110110,
        48'b110110110110110110110110110110110110110110110110,
        48'b110110110110110110110110110110110110110110110110,
        //tile_code 63
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010001010011010010010010010010010011010010001011,
        48'b011001001001001001001001001001001001001001001011,
        48'b010001100100100100100100011011010010100100001011,
        48'b010001100100100100011010010010011011011100001011,
        48'b010001100100100010010011010011011011101110001011,
        48'b011001100100010011010010011011100101101110001011,
        48'b010001100010010010011011011100100011010010001011,
        48'b010001010010010011011101101110110010011011001011,
        48'b010001011011011100101101101011010010011100001011,
        48'b011001101110100100110011010010011011100100001011,
        48'b010001100110110010010010011011100100100100001011,
        48'b010001001001001001001001001001001001001001001011,
        48'b000001000000000000000000000000000000000000001000,
        48'b001001001001001001001001001001001001001001001001,
        //tile_code 64
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001010010001001010010001001010010001001000,
        48'b000001001010010001001010010001001010010001001000,
        48'b000001001010010001001010010001001010010001001000,
        48'b000011000100100011000100100011000100100011000000,
        48'b000000011011011000011011011000011011011000011000,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b101110101111111111111111111101110110110110110101,
        48'b101110101111111111111111111101110101101101110101,
        48'b101110101111111111111111111101110101111101110101,
        48'b101110101111111111111111111101110101111101110101,
        48'b101110101111111111111111111101110101101101110101,
        48'b101110101111111111111111111101110111111111110101,
        48'b101110101111111111111111111101110101101101110101,
        48'b101110101111111111111111111101110101111101110101,
        //tile_code 65
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010001010010010010010010010010010010010010001010,
        48'b011001001001001001001001001001001001001001001011,
        48'b010001100100100100100100101101101101100100001010,
        48'b010001100100100100100110101101101101101100001010,
        48'b010001100100100100100110110110101101101100001010,
        48'b011001100100100100110101110110110110111100001011,
        48'b010001100100100110110110110101111111101100001010,
        48'b010001100100100110101110111111111101101100001010,
        48'b010001100100110110111111111101101111101100001010,
        48'b011001100110111111111101101111101101100100001011,
        48'b010001100111111101101111101101100100100100001010,
        48'b010001001001001001001001001001001001001001001010,
        48'b000001000000000000000000000000000000000000001000,
        48'b001001001001001001001001001001001001001001001001,
        //tile_code 66
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        //tile_code 67
        48'b000000001001001001001001001010010010010010000000,
        48'b000000001001001001001001001000000000000000000000,
        48'b000000001001001001001001001001001001001011000000,
        48'b000000001001001001001001001001001001011011000000,
        48'b000000001001001001001001001001001011011001000000,
        48'b000000001001001001001001001001011011001001000000,
        48'b000000001001001001001001001011011001001001000000,
        48'b000000001001001001001001011011001001001011000000,
        48'b000000001001001001001011011001001001011001000000,
        48'b000000001001001001011011001001001011001001000000,
        48'b000000001001001011011001001001011001001001000000,
        48'b000000001001011011001001001011001001001001000000,
        48'b000000010011011010010010011010010010010010000000,
        48'b000000011011010010010011010010010010010010000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 68
        48'b000000001001001001001010010010010010010010000000,
        48'b000000000000000000000010010010010010010010000000,
        48'b000000010010010010010010010010010010010011000000,
        48'b000000010010010010010010010010010010011011000000,
        48'b000000010010010010010010010010010011011010000000,
        48'b000000010010010010010010010010011011010010000000,
        48'b000000010010010010010010010011011010010010000000,
        48'b000000010010010010010010011011010010010011000000,
        48'b000000010010010010010011011010010010011010000000,
        48'b000000010010010010011011010010010011010010000000,
        48'b000000010010010011011010010010011010010010000000,
        48'b000000010010011011010010010011010010010010000000,
        48'b000000001011011001001001011001001001001001000000,
        48'b000000011011001001001011001001001001001001000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 69
        48'b000001001001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010010010010010010010010010010010010010010,
        48'b000010010010010010010010010010010010010010010010,
        48'b000001001001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010010010010010010010010010010010010010010,
        48'b000010010010010010010010010010010010010010010010,
        48'b000001001001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010010010010010010010010010010010010010010,
        48'b000010010010010010010010010010010010010010010010,
        48'b000001001001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010010010010010010010010010010010010010010,
        48'b000010010010010010010010010010010010010010010010,
        //tile_code 70
        48'b000001010010010010010010010010010011100100011000,
        48'b000001000000000000000000000000000011011011011000,
        48'b000001000101101101101101101101101011100100011000,
        48'b000001000001001001001001001001001011110110011000,
        48'b000001000001001001001001001001001001011011001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000000000000000000000000000000000000001000,
        48'b000001000000000000000000000000000000000000001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 71
        48'b000001001001001001001001001001001001001001001000,
        48'b000010010001010010010010010010010010010010010000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000010010010010010010010010010010001010010010000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000010010010010001010010010010010010010010010000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000010010010010010010010010010001010010010010000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 72
        48'b000001001001001001001001001001001001001001001001,
        48'b001010001011011011011011011011011011011011011011,
        48'b001001001000000000000000000000000000000000000000,
        48'b001000001100100100100100100100100100100100100100,
        48'b001000001100100100100100100100100100100100100100,
        48'b001001001000000000000000000000000000000000000000,
        48'b001101001110110110110110110110110110110110110110,
        48'b001101001100100100100100100100100100100100100100,
        48'b001101001110110110110110110110110110110110110110,
        48'b001001001000000000000000000000000000000000000000,
        48'b001000001100100100100100100100100100100100100100,
        48'b001001001001001001001001001001001001001001001001,
        48'b001000000001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b010010010010010010010000010010010010010010010000,
        48'b101101101101101101101101101101101101101101101101,
        //tile_code 73
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010000011000,
        48'b001001001001001001001001001001001001001000000000,
        48'b100100100100100100100100100100100100100000001000,
        48'b100100100100100100100100100100100100100000001000,
        48'b001001001001001001001001001001001001001000000000,
        48'b101101101101101101101101101101101101101000110000,
        48'b100100100100100100100100100100100100100000110000,
        48'b101101101101101101101101101101101101101000110000,
        48'b001001001001001001001001001001001001001000000000,
        48'b100100100100100100100100100100100100100000001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000000000001,
        48'b011011011011011011011001011011011011011011011001,
        48'b110110110110110110110110110110110110110110110110,
        //tile_code 74
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000010010010010000001000000000000,
        48'b011011011011011010100100100100010011011011011011,
        48'b000000000000010101110110110110101010000000000001,
        48'b000000000000001010101101101101010001000000000001,
        48'b000000000000010001010010010010001010000000000001,
        48'b011011011011010010010010010010010010011011011011,
        48'b000000000001010001011001001011001010000000000000,
        48'b000000000001010001011001001011001010000000000000,
        48'b000000000001010001011001001011001010000000000000,
        48'b011011011011011010001001001001010011011011011011,
        48'b000000000000000000010010010010000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b011011011011011011011011011011011011011011011011,
        //tile_code 75
        48'b000001001000001001001001001001001000001001001000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000011011011011011011011011011011011011011011000,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011000,
        48'b000001001000001001001001001001001000001001001000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000011011011011011011011011011011011011011011000,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011000,
        //tile_code 76
        48'b000001000010010010010010010000001000010000001000,
        48'b000001000010010010010010010000001000000000001000,
        48'b000001000010010010010010010000001000010000001000,
        48'b000001000010010010010010010000001000000000001000,
        48'b000001000010010010010010010000001000000000001000,
        48'b000001000010010010010010010000001000000000001000,
        48'b000001000000000000000000000000001000000000001000,
        48'b000001000000000000000000000000001000010000001000,
        48'b000001001001001001001001001001001000000000001000,
        48'b000001000000000000000000000000001010010010001000,
        48'b000001000010010010010010010000001001001001001000,
        48'b000001000010010010010010010000001001001001001000,
        48'b000001000000000000000000000000001001001001001000,
        48'b000001000000000000000000000000001001001001001000,
        48'b000010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 77
        48'b000001000010000001000010010010010010010000001000,
        48'b000001000000000001000010010010010010010000001000,
        48'b000001000010000001000010010010010010010000001000,
        48'b000001000000000001000010010010010010010000001000,
        48'b000001000000000001000010010010010010010000001000,
        48'b000001000000000001000010010010010010010000001000,
        48'b000001000000000001000000000000000000000000001000,
        48'b000001000010000001000000000000000000000000001000,
        48'b000001000000000001001001001001001001001001001000,
        48'b000001010010010001000000000000000000000000001000,
        48'b000001001001001001000010010010010010010000001000,
        48'b000001001001001001000010010010010010010000001000,
        48'b000001001001001001000000000000000000000000001000,
        48'b000001001001001001000000000000000000000000001000,
        48'b000010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 78
        48'b000000000001000000010010010010000001000000000000,
        48'b000000000010010010011011011011010010010000000000,
        48'b000000010011011100101101101101100011011010000000,
        48'b110010011101101111100100100100111101101011010110,
        48'b010111100101101100101101101101100101101100111010,
        48'b010111101100100100111111111111100100100101111010,
        48'b000010101101101111100100100100111101101101010001,
        48'b010111100111111100101101101101100111111100111010,
        48'b010111101100100100111111111111100100100101111010,
        48'b000010101101101111100100100100111101101101010000,
        48'b000000010111111100111101101111100111111010000000,
        48'b110010111100100100111111111111100100100111010110,
        48'b010010111111111111100100100100111111111111010010,
        48'b010010010111111100111111111111100111111010010010,
        48'b010010010010010010111111111111010010010010010010,
        48'b110010010010010010010010010010010010010010010110,
        //tile_code 79
        48'b000001001001001001001001001001001001001001001010,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000010010010010010010010010010010010010010010010,
        48'b011000000000000000000000000000000000000000000000,
        //tile_code 80
        48'b000001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b000000000000000000000000000000000000000000000010,
        48'b010010010010010010010010010010010010010010010011,
        //tile_code 81
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000010010010010010010010010010010010010010010000,
        48'b011000000000000000000000000000000000000000000000,
        //tile_code 82
        48'b000001001001001001001001001001001001001001001010,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000010010010010010010010010010010010010010010011,
        48'b000010011011011011011011011011011011011011010011,
        //tile_code 83
        48'b000001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b000000000000000000000000000000000000000000000010,
        48'b011000011011011011011011011011011011011011000010,
        //tile_code 84
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000011011011011011011011011011011011011011011011,
        48'b011100100100100100100101101101101101101101101101,
        48'b011100100011011011011011011011011011011011011100,
        48'b011100100011011011011011011011011011011011011100,
        48'b011100011101101101101101101101101101101101101100,
        48'b011100011101101101101101101101101101101101101100,
        48'b011100011101101101101101101101101101101101101100,
        48'b011101011101110110110110110110110110110110110100,
        48'b011101011101110110110110110110110110110110110100,
        48'b011101011101110110110110110110110110110110110100,
        48'b011101011101110110110110110110110110110110110100,
        //tile_code 85
        48'b000000000001001001001001001001001001001001001001,
        48'b000000001010010010010010010010010010010010010010,
        48'b000001010010011011011011011011011011011011011011,
        48'b001010100010011011011011011011011011011011011011,
        48'b001010100010011011011011011011011011011011011011,
        48'b010100100010011011011011011011011011011011011011,
        48'b100100100010011011011011011011011011011011011011,
        48'b100100100010011011011011011011011011011011011011,
        48'b100100100010011011011011011011011011011011011011,
        48'b100100100010011011011011011011011011011011011011,
        48'b100100100010011011011011011011011011011011011011,
        48'b100100100010011011011011011011011011011011011011,
        48'b100100100010011011011011011011011011011011011011,
        48'b100100100010010011011011011011011011011011011011,
        48'b100100100010010011011011011011011011011011011011,
        48'b100100101001001001001001001001001001001001001001,
        //tile_code 86
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 87
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 88
        48'b000000000001000000000000000000010010000000000000,
        48'b000000000001000000000000000010011011010000000000,
        48'b000000000001000000000000010011100100011010010000,
        48'b101101101101101101010010010011100100011010110010,
        48'b000000000000000010110110010011010010011010111010,
        48'b000000000000000010111111111010111010010010010001,
        48'b000000000000000000010010010010010000000000000001,
        48'b101101101101101101101101101101101101101101101101,
        48'b000000000001000010010000000000000001000000000000,
        48'b000000000001010011011010000000000001000000000000,
        48'b000000000010011100100011010010000001000000000000,
        48'b101010010010011100100011010110010101101101101101,
        48'b010110110010011010010011010111010000000000000001,
        48'b010111111111010111010010010010000000000000000001,
        48'b000010010010010010000001000000000000000000000001,
        48'b101101101101101101101101101101101101101101101101,
        //tile_code 89
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000011011000000000000001,
        48'b000000000000000000000001000011000000000000000001,
        48'b010010010010010010010010010011000011010010010010,
        //tile_code 90
        48'b000001000001010010010010010010010010010010010011,
        48'b000001000001010010010010010010010010010010010011,
        48'b000001000001010010010010010010010010010010010011,
        48'b000001000001001001001010010010010010010010010011,
        48'b000000000000000000000000000000000000000000000000,
        48'b000011011011011011011011011011011011011011011011,
        48'b000010010010010010010010010010010010010010010010,
        48'b000010010010010010010010010010010010010010010010,
        48'b000010010010010010010000000000000000000000000000,
        48'b000010010010010010010000000000000000000000000000,
        48'b100000000000000000000000011010010010010010010001,
        48'b101000010010010010000000000000000000000000000000,
        48'b100100000000000000000110110110100110100110100110,
        48'b100100110110110110110000000111111111111111111000,
        48'b100100110110110110110000000111111111111111111000,
        48'b101101101110110110110110110000000000000000000110,
        //tile_code 91
        48'b000001010010010010010010010010010010010010010010,
        48'b001010001011011010000000000000000000000000000010,
        48'b010100100011011010000000000000000000000000000010,
        48'b010100100011011010000000000000000000000000000010,
        48'b001011011011010010010010010010010010010010010011,
        48'b001100100011010001001001001001001001010010001011,
        48'b100100100011010001101101101101101101101101101011,
        48'b100100100011010001001001101101101101101101101011,
        48'b011100100011010001001001101101101101101101101011,
        48'b011100100011010001001001101101101101101101101011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011100100100100100100100100100100100100100100,
        48'b110011011011011011011011011011011011011011011011,
        48'b011110110110110110110110110110110110110110110110,
        48'b011110110110110110110110110110110110110110110110,
        48'b110110110110110110110110110110110110110110110110,
        //tile_code 92
        48'b000000000000000000000000000000000000000000000000,
        48'b001010010010010010010010010010010010010010010010,
        48'b001010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010011011,
        48'b010010010010010010010010010010010010010010011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b010010010010010010010010010010010010010010011011,
        48'b011011011011011011011011011011011011011011011100,
        48'b101101101101101101101101101101101101101101101011,
        48'b101101101101101101101101101101101101101101101011,
        48'b101101101101101101101101101101101101101101101101,
        //tile_code 93
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b001001001001001001001001001010010010010010010001,
        48'b001001001001001001001001001010010010010010010001,
        48'b000010010010010010010000001001001001001001001001,
        48'b001001001001001001001001001001010010010010001011,
        48'b100100011100011100011100100001001001001001100101,
        48'b001101101101101101101001001100100100100100100101,
        48'b001101101101101101101001001100100100100100100101,
        48'b100001001001001001001100100100100100100100011011,
        //tile_code 94
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000010010000000001000000000000,
        48'b000000000001000000010000000010000001000000000000,
        48'b011011011011011011010000000010011011011011011011,
        48'b000000000000000000010000000010000000000000000001,
        48'b000000000000000010000000000000010000000000000001,
        48'b000000000000000010000000000000010000000000000001,
        48'b011011011011011010011011011011010011011011011011,
        48'b000000000001000100010010010010100001000000000000,
        48'b000000000001000100101110110101100001000000000000,
        48'b000000000001000000100100100100000001000000000000,
        48'b011011011011011011010011011010011011011011011011,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b011011011011011011010011011010011011011011011011,
        //tile_code 95
        48'b000000000001000000000000000010000011010000000000,
        48'b000000000001000000000010010010010001010000000000,
        48'b000000000001000000010000000010010010000000000000,
        48'b011011011011011011010000000010010011010011011011,
        48'b000000000000000000010000000010010001010000000001,
        48'b000000000000000000010000000010010010000000000001,
        48'b000000000000000000010001001010010011010000000001,
        48'b011011011011011011010011011010010001010011011011,
        48'b000000000001000000001010010010010010000000000000,
        48'b000000000001000000010011011010010001000000000000,
        48'b000000000001000000010011011010010001000000000000,
        48'b011011011011011011010011011010011011011011011011,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b011011011011011011010011011010011011011011011011,
        //tile_code 96
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000011011000000000000000000001,
        48'b010010010010010010011010010011010010010010010010,
        48'b000000000001000000011010010011000001000000000000,
        48'b000000000001000000001011011001000001000000000000,
        48'b000000000001000000011001001011000001000000000000,
        48'b010010010010010010010011011010010010010010010010,
        48'b000000000000000000011000000011000000000000000001,
        48'b000000000000000000011011011011000000000000000001,
        48'b000000000000000000011001001011000000000000000001,
        48'b010010010010010010011001001011010010010010010010,
        //tile_code 97
        48'b000000000001000000000010010000000001000000000000,
        48'b000000000001000000010000000010000001000000000000,
        48'b000000000001000000010000000010000001000000000000,
        48'b011011011011011011010000000010011011011011011011,
        48'b000000000000000010000000000000010000000000000001,
        48'b000000000000000010000000000000010000000000000001,
        48'b000000000000000010011011011011010000000000000001,
        48'b011011011011011100010010010010100011011011011011,
        48'b000000000001000100101110110101100001000000000000,
        48'b000000000001000000100100100100000001000000000000,
        48'b000000000001000000010011011010000001000000000000,
        48'b011011011011011011010011011010011011011011011011,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b011011011011011011010011011010011011011011011011,
        //tile_code 98
        48'b000000000001000000010011011010000001000000000000,
        48'b000000000001000000010011011010000001000000000000,
        48'b000000000001000000010011011010000001000000000000,
        48'b011011011011011011010011011010011011011011011011,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b011011011011011011010011011010011011011011011011,
        48'b000000000001000000010011011010000001000000000000,
        48'b000000000001000000010011011010000001000000000000,
        48'b000000000001000000010011011010000001000000000000,
        48'b011011011011011011010011011010011011011011011011,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b011011011011011011010011011010011011011011011011,
        //tile_code 99
        48'b000000000001000000010011011010000001000000000000,
        48'b000000000001000000011000000011000001000000000000,
        48'b000000000001000000011011011011000001000000000000,
        48'b010010010010010010011001001011010010010010010010,
        48'b000000000000000000011001001011000000000000000001,
        48'b000000000000000000011001001011000000000000000001,
        48'b000000000000000000011001001011000000000000000001,
        48'b010010010010010010011001001011010010010010010010,
        48'b000000000001000000011001001011000001000000000000,
        48'b000000000001000000011001001011000001000000000000,
        48'b000000000001000000001011011001000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        //tile_code 100
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000010010000000001000000000000,
        48'b011011011011011011011010010011011011011011011011,
        48'b000000000000000000000010010000000000000000000001,
        48'b000000000000000000010100100010000000000000000001,
        48'b000000000000000000010101101010000000000000000001,
        48'b011011011011011011010101101010011011011011011011,
        48'b000000000001010010100100100100010010000000000000,
        48'b000000000010100010101100100101010100010000000000,
        48'b000000000010100010101101101101010100010000000000,
        48'b011011011010110110100101101100110110010011011011,
        48'b000000000111010010110110110110010010111000000001,
        48'b000000000000111111010010010010111111000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b011011011011011011011011011011011011011011011011,
        //tile_code 101
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000010010010010000001000000000000,
        48'b011011011011010010100100100100010010011011011011,
        48'b000000000010100100010010010010100100010000000001,
        48'b000000000010100010010100010100010100010000000001,
        48'b000000010100010010100010100010100010100010000001,
        48'b011011010100010100010100010100010010100010011011,
        48'b000000010100010010100010100010100010100010000000,
        48'b000000000010100010010100010100010100010000000000,
        48'b000000000010100100010010010010100100010000000000,
        48'b011011011011010010100100100100010010011011011011,
        48'b000000000000000000010010010010000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b011011011011011011011011011011011011011011011011,
        //tile_code 102
        48'b000000000000000000000001001000000000000000000000,
        48'b000010010010010010000001001000010010010010010001,
        48'b000010010010010010000001001000010010010010010011,
        48'b000010010010010010000001001000010010010010010011,
        48'b000010010010010010000001001000010010010010010011,
        48'b000010010010010010000001001000010010010010010000,
        48'b000010010010010000000001001000000010010010010000,
        48'b000010010010000001000001001000001000010010010000,
        48'b000010010000001001011001001011001001000010010000,
        48'b000010010010000011011011011011011000010010010000,
        48'b000010010010010000000000000000000010010010010000,
        48'b000010010010010010000000000000010010010010010000,
        48'b000010010010010010000000000000010010010010010000,
        48'b000010010010010010000000000000010010010010010000,
        48'b000001001001001001000000000000001001001001001000,
        48'b000001011011011011000000000000011011011011001000,
        //tile_code 103
        48'b000000000000000000000001001000000000000000000000,
        48'b010010010010010010000001001000010010010010010001,
        48'b010010010010010010000001001000010010010010010011,
        48'b010010010010010010000001001000010010010010010011,
        48'b010010010010010010000001001000010010010010010011,
        48'b010010010010010010000001001000010010010010010011,
        48'b010010010010010000000001001000000010010010010011,
        48'b010010010010000001000001001000001000010010010011,
        48'b010010010000001001011001001011001001000010010011,
        48'b010010010010000011011011011011011000010010010011,
        48'b010010010010010000000000000000000010010010010011,
        48'b010010010010010010000000000000010010010010010011,
        48'b010010010010010010000000000000010010010010010011,
        48'b010010010010010010000000000000010010010010010011,
        48'b001001001001001001000000000000001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 104
        48'b000000000000000000000001001000000000000000000000,
        48'b010010010010010010000001001000010010010010010001,
        48'b010010010010010010000001001000010010010010010011,
        48'b010010010010010010000001001000010010010010010011,
        48'b010010010010010010000001001000010010010010010011,
        48'b010010010010010000000001001000000010010010010011,
        48'b010010010010000001000001001000001000010010010011,
        48'b010010010000001001011001001011001001000010010011,
        48'b010010010010000011011011011011011000010010010011,
        48'b010010010010010000000000000000000010010010010011,
        48'b010010010010010010000000000000010010010010010011,
        48'b010010010010010010000000000000010010010010010011,
        48'b010010010010010010000000000000010010010010010011,
        48'b010010010010010010000000000000010010010010010011,
        48'b001001001001001001000000000000001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 105
        48'b000000000000000000000001001000000000000000000000,
        48'b010010010010010010000001001000010010010010010000,
        48'b010010010010010010000001001000010010010010010000,
        48'b010010010010010010000001001000010010010010010000,
        48'b010010010010010010000001001000010010010010010000,
        48'b010010010010010000000001001000000010010010010000,
        48'b010010010010000001000001001000001000010010010000,
        48'b010010010000001001011001001011001001000010010000,
        48'b010010010010000011011011011011011000010010010000,
        48'b010010010010010000000000000000000010010010010000,
        48'b010010010010010010000000000000010010010010010000,
        48'b010010010010010010000000000000010010010010010000,
        48'b010010010010010010000000000000010010010010010000,
        48'b010010010010010010000000000000010010010010010000,
        48'b001001001001001001000000000000001001001001001000,
        48'b000001011011011011000000000000011011011011001000,
        //tile_code 106
        48'b000000000000000000000001001000000000000000000000,
        48'b000010010010010010000001001000010010010010010001,
        48'b000010010010010010000001001000010010010010010011,
        48'b000010010010010010000001001000010010010010010011,
        48'b000010010010010010000001001000010010010010010011,
        48'b000010010010010010000001001000010010010010010011,
        48'b000010010010010000000001001000000010010010010011,
        48'b000010010010000001000001001000001000010010010011,
        48'b000010010000001001011001001011001001000010010011,
        48'b000010010010000011011011011011011000010010010011,
        48'b000010010010010000000000000000000010010010010011,
        48'b000010010010010010000000000000010010010010010011,
        48'b000010010010010010000000000000010010010010010011,
        48'b000010010010010010000000000000010010010010010011,
        48'b000001001001001001000000000000001001001001001001,
        48'b000001011011011011000000000000011011011011001000,
        //tile_code 107
        48'b000001001001001001000000000000001001001001001010,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000010001001001001000000000000001001001001001011,
        48'b011000001001001001001000000001001001001001001011,
        48'b011000010001001001001001001001001001001001001011,
        48'b011011000010010001001001001001001001001001001011,
        48'b011011011000000010010010010010010010010010010010,
        48'b011011011011011000000000000000000000000000000000,
        //tile_code 108
        48'b000001010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010001,
        48'b010010010010010010000000000000010010010010010000,
        48'b010010010010010010000000000000010010010010001000,
        48'b010010010010010010000000000000010010001001000011,
        48'b001001001001001001000000000000001001000000011011,
        48'b000000000000000000000000000000000000011011011011,
        //tile_code 109
        48'b000001001001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b000001010010010010010010010010010010010010010010,
        48'b000001010010010010010010010010010010010010010010,
        48'b000001010010001001001001001001001001001001001001,
        48'b000001010010001001001001001001001001001001001001,
        48'b000001010010001001001001001001001001001001001001,
        48'b000001010010001001001001001001001001001001001001,
        48'b000001010010001001001001001001001001001001001001,
        48'b000001010010001001001001001001001001001001001001,
        48'b000001010010001001001001001001001001001001001001,
        48'b001001010010001001001001001001001001001001001001,
        48'b001001010010010010001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001010010010010010010010010001001001001,
        //tile_code 110
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile_code 111
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001001001000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile_code 112
        48'b000000000000000000001001001001000000000000000000,
        48'b000000000000000000001001001001000000000000000000,
        48'b010010010010010010001001001001010010010010010010,
        48'b010010010010010010001001001001010010010010010010,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000000001001000000000000000000000,
        48'b010010010000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000010010010010010010010010000000000000,
        //tile_code 113
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile_code 114
        48'b000000000000000000001001001001000000000000000000,
        48'b000000000000000000001001001001000000000000000000,
        48'b010010010010010010001001001001010010010010010010,
        48'b010010010010010010001001001001010010010010010010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000000001001000000000000000000010,
        48'b000000000000000000000000000000000000000010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000010010010010010010010010000000000000,
        //tile_code 115
        48'b000000000000000000001001001001000000000000000000,
        48'b000000000000000000001001001001000000000000000000,
        48'b010010010010010010001001001001010010010010010010,
        48'b010010010010010010001001001001010010010010010010,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000000001001000000000000000000000,
        48'b010000000000000000000000000000000000000000000000,
        48'b010010010000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000010010010010010010010010000000000000,
        //tile_code 116
        48'b000000000000000000001001001001000000000000000000,
        48'b000000000000000000001001001001000000000000000000,
        48'b010010010010010010001001001001010010010010010010,
        48'b010010010010010010001001001001010010010010010010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000000001001000000000000000000010,
        48'b000000000000000000000000000000000000000000000010,
        48'b000000000000000000000000000000000000000010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000010010010010010010010010000000000000,
        //tile_code 117
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001000,
        48'b001001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile_code 118
        48'b000001001001001001000000000000001001001001001010,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000010001001001001001000000001001001001001001011,
        48'b011000001001001001001001001001001001001001001011,
        48'b011000010001001001001001001001001001001001001011,
        48'b011011000010010001001001001001001001001001001011,
        48'b011011011000000010010010010010010010010010010010,
        48'b011011011011011000000000000000000000000000000000,
        //tile_code 119
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile_code 120
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        //tile_code 121
        48'b000000000000000000001001001001000000000000000000,
        48'b000000000000010010001001001001010010000000000000,
        48'b000000000000010010001001001001010010000000000000,
        48'b000000000000010010001001001001000000000000000000,
        48'b000000000000010010001001001001000000000000000000,
        48'b000000000000010010000001001000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010010010010010010010000000000000,
        //tile_code 122
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile_code 123
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b010010010010010010010010010010001001000000000000,
        48'b010010010010010010010010010010001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        //tile_code 124
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001010010010010010010010010010010,
        48'b000000000000001001010010010010010010010010010010,
        48'b000000000000001001000000000000000000000000000000,
        //tile_code 125
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 126
        48'b000000000000000000000000000000001001000000000000,
        48'b010010010010010010010010010010001001000000000000,
        48'b010010010010010010010010010010001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile_code 127
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001010010010010010010010010010010,
        48'b000000000000001001010010010010010010010010010010,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile_code 128
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000010010010010010010010010000000000000,
        //tile_code 129
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 130
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 131
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 132
        48'b000000000000000001001001001001001001001001001001,
        48'b000000000001001010010010010010010010010010010011,
        48'b000000001010010010010010010010010010010010010000,
        48'b000001010010010010010010010010010010010010010000,
        48'b000001010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001011011011011011011011011011011011011011011000,
        48'b001011000000000000000000000000000000000000000011,
        //tile_code 133
        48'b000000000000000000000000000000000001001001001001,
        48'b010010010010010010010010010010010000000001001001,
        48'b010010010010010010010010010010010010010000001001,
        48'b010010010010010010010010010010010010010010000001,
        48'b010010010010010010010010010010010010010010000001,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011001001001001001001001001001001001001001011000,
        //tile_code 134
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 135
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000001001001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 136
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 137
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000001001001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b001001001001001001001001001001001001001001001000,
        48'b001001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 138
        48'b000001001001001001001001001001001001001001001000,
        48'b010001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b010010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 139
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001010,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001000000001001001001011,
        48'b000010010010010010010010010000001010010010010010,
        48'b000000000000000000000000000000001000000000000000,
        //tile_code 140
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b010010010010010010010010010010010010010010010010,
        48'b011000000000000000000000000000000000000000000000,
        //tile_code 141
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000011,
        //tile_code 142
        48'b000001001001001001001001001001001001001001001001,
        48'b001010010010010010010010010010010010010010010011,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001011011011011011011011011011011011011011011000,
        48'b001011000000000000000000000000000000000000000011,
        //tile_code 143
        48'b000001001001001001001001001001001001001001001001,
        48'b001010010010010010010010010010010010010010010011,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010001001010010010010000,
        48'b001011011011011011011011011001010011011011011000,
        48'b001011000000000000000000000001010001000000000011,
        //tile_code 144
        48'b000001000010010010010010010010010010010010010010,
        48'b000000000011011011011011011011011011011011011011,
        48'b000011000100100100100100100100100100100100100100,
        48'b000011000100100100100100100100100100100100100100,
        48'b000000000011011011011011011011011011011011011011,
        48'b000101000110110110110110110110110110110110110110,
        48'b000101000100100100100100100100100100100100100100,
        48'b000101000110110110110110110110110110110110110110,
        48'b000000000011011011011011011011011011011011011011,
        48'b000011000100100100100100100100100100100100100100,
        48'b000000000000000000000000000000000000000000000000,
        48'b000011011000000000000000000000000000000000000000,
        48'b011000000000000000000000000000000000000000000000,
        48'b001001001001001001001011001001001001001001001011,
        48'b001001001001001001001011001001001001001001001011,
        48'b101101101101101101101101101101101101101101101101,
        //tile_code 145
        48'b000000000000000000000000000000000000000001010001,
        48'b011011011011011011011011011011011011011001001001,
        48'b100100100100100100100100100100100100100001011001,
        48'b100100100100100100100100100100100100100001011001,
        48'b011011011011011011011011011011011011011001001001,
        48'b101101101101101101101101101101101101101001110001,
        48'b100100100100100100100100100100100100100001110001,
        48'b101101101101101101101101101101101101101001110001,
        48'b011011011011011011011011011011011011011001001001,
        48'b100100100100100100100100100100100100100001011001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001011011001,
        48'b001001001001001001001001001001001001001001001011,
        48'b010010010010010010010011010010010010010010010011,
        48'b010010010010010010010011010010010010010010010011,
        48'b110110110110110110110110110110110110110110110110,
        //tile_code 146
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001010010001001001001001001001,
        48'b001001001001001001001010010001001001001001001001,
        48'b001000000000000000000010010000000000000000000000,
        48'b001000000000000000010011011010000000000000000000,
        48'b001000000000000000010001001010000000000000000000,
        48'b001000000000000000010001001010000000000000000000,
        48'b001000000000010010011011011011010010000000000000,
        48'b001000000010011010001011011001010011010000000000,
        48'b001000000010011010001001001001010011010000000000,
        48'b001000000010100100011001001011100100010000000000,
        48'b001001001101010010100100100100010010101000000000,
        48'b000000000000101101010010010010101101000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile_code 147
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001010,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 148
        48'b000001001001001001001001001001001001001001001001,
        48'b001010011011011011011011011011011011011011011011,
        48'b001010010010010010010010010010010010010010010010,
        48'b001010010000001001001001001001001001001001001001,
        48'b001010010001100100100100100100100100100100100100,
        48'b001010010001100100100100100100100100100100100100,
        48'b001010010001100100100100100100100100100100100100,
        48'b001010010001100100100100100100100100100100100100,
        48'b001010010001100100100100100100100100100100100100,
        48'b001010010001100100100100100100100100100100100100,
        48'b001010010001001001001001001001001001001001001001,
        48'b001010010001010010010010010010010010010010010010,
        48'b001010010001010010010010010010010010010010010010,
        48'b001010010001010010010010010010010010010010010010,
        48'b001010010001010010010010010010010010010010010010,
        48'b001010010001010010010010010010010010010010010010,
        //tile_code 149
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        //tile_code 150
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010000,
        48'b011011011011011011011011011011011011011011011000,
        48'b000000000000000000000000000000000000001011011000,
        48'b100100100100100100100100100100100100000011011000,
        48'b100100100100100100100100100100100100000011011000,
        48'b100100100100100100100100100100100100000011011000,
        48'b100100100100100100100100100100100100000011011000,
        48'b100100100100100100100100100100100100000011011000,
        48'b100100100100100100100100100100100100000011011000,
        48'b000000000000000000000000000000000000000011011000,
        48'b011011011011011011011011011011011011000011011000,
        48'b011011011011011011011011011011011011000011011000,
        48'b011011011011011011011011011011011011000011011000,
        48'b011011011011011011011011011011011011000011011000,
        48'b011011011011011011011011011011011011000011011000,
        //tile_code 151
        48'b000001001000000001001000000001001000000001001000,
        48'b001010011001001010011001001010011001001010011001,
        48'b001001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b001010011000000010011000000010011000000010011000,
        48'b001010011000000010011000000010011000000010011000,
        48'b001001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b001010011000000010011000000010011000000010011000,
        48'b001010011000000010011000000010011000000010011000,
        48'b001001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b001010011000000010011000000010011000000010011000,
        48'b001010011000000010011000000010011000000010011000,
        48'b001001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        //tile_code 152
        48'b000001001000000001001000000001001000000001001000,
        48'b001010011001001010011001001010011001001010011001,
        48'b000001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011000,
        48'b000010011000000010011000000010011000000010011000,
        48'b000001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011000,
        48'b000010011000000010011000000010011000000010011000,
        48'b000001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011000,
        48'b000010011000000010011000000010011000000010011000,
        48'b000001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        //tile_code 153
        48'b000001001000000001001000000001001000000001001000,
        48'b001010011001001010011001001010011001001010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001000000001001000000001001000000001001000000001,
        //tile_code 154
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000011000000001000000000000000000000001,
        48'b010010010011011011010010010010010010010010010010,
        48'b000000000001011000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000100100100000000000000,
        48'b010010010010010010010100100100100100100100100101,
        48'b000000000000000000100100100100110110110110100011,
        48'b000000000000100100100110110111110110100011101101,
        48'b000000000100100100110111111111110111011101101101,
        48'b100100100100111111110111111111110110110110101101,
        //tile_code 155
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000011011011011011000000000000000001000000000000,
        48'b011011011011011100100100100100100100010010010010,
        48'b100011011011101100100100100100100100100011011011,
        48'b100101101101101101101101100100100100100011011011,
        48'b100100101101101101101101101101100100100100011011,
        48'b100100100101101101101101101101101101101100011011,
        //tile_code 156
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010011010010010010010010010010010,
        48'b000000000001000011011011000000000001000000000000,
        48'b000000000001000000011000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b100000000000000000000001000000000000000000000001,
        48'b100100100100100100100100100000000000000000000001,
        48'b100100100100100100100100100100100100100000101101,
        48'b100100100100011101101101101101101100101101101101,
        //tile_code 157
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010011011011011011010010010010010010,
        48'b000000000000011011011011011011011000000000000001,
        48'b000000000000000011011011011011000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b100100100100100000000101101101101101101101101001,
        48'b100100100100100101101101101101101101101101101101,
        //tile_code 158
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000011,
        48'b000000000001000000000000000000000001000000011011,
        48'b000000000001000000000000000000000011011011011011,
        48'b010010010010010010010010010010011011011011011011,
        48'b000000000000000000000001000011011011011011011011,
        48'b000000000000000000000001000000011011011011011011,
        48'b000000000000000000000001000000000000011011011011,
        48'b100100100010010010010010010010010010010010010010,
        //tile_code 159
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011000001000000000000000000000001000000000000,
        48'b011011011001000000000000000000000001000000000000,
        48'b011011011011000000000000000000000001000000000000,
        48'b011011011010010010010010010010010010010010010100,
        48'b011011000000000000000001000100100100100100100100,
        48'b011000000000000000000100100100100100100100100100,
        48'b000000000000000000100100100100100100100100100100,
        48'b010010010010010100100100100100100100100100100100,
        //tile_code 160
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000011011011,
        48'b010010010010010010010010010010010011011011011011,
        48'b000000000001000000000000000011011011011011011011,
        48'b000000000001000000000000000011011011011011011011,
        48'b100100100100100100100000000011011011011011011011,
        48'b100100100100100100100100011011011011011011011011,
        48'b100100100100100100100011011011011011011011011011,
        48'b100100100100100100011011011011011011011011011011,
        48'b100100100100011011011011011101011011011011011011,
        48'b100100011011011011011101101101101011011011011011,
        //tile_code 161
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b011011000000000000000001000000000000000000000001,
        48'b011011011010010010010010010010010010010010010010,
        48'b011011011011011011000000000000000001000000000000,
        48'b011011011011011011011011011000000001011011011000,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011100011100011011011011011011011011011,
        48'b011011011100100100100100011011011011011011011011,
        //tile_code 162
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000011011011011000000000000000001000000000000,
        48'b100011011011011011011010010010010010010010010010,
        48'b100100011011011011011011000000000000000000000001,
        48'b100100011011101011011011011000000000000000011011,
        48'b100100100110101011100100100000000000000011011011,
        48'b100100110101101100100100100100100011011011011011,
        //tile_code 163
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000011000000000001000000000000000000000001,
        48'b000000011011011011011011000000000000000000000001,
        48'b010010011011011011011011011010010010010010010010,
        48'b000000000011011011011011000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000100100100100100100100100100100100100000001,
        48'b100100100100100100100100100100100100100100100100,
        48'b100100100100100100100100100100100100100100100100,
        48'b100100100100100100100100100100100100100100100100,
        //tile_code 164
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b011011000000000000000001000000000000000000000001,
        48'b011011011011011000100100100100100100100100100100,
        48'b011011011011100100100100100100100100100100100100,
        //tile_code 165
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b011011011000000000000001000000000000000000000001,
        48'b011011011011011011011011010010010010010010010010,
        //tile_code 166
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010011011011011011011011011011010010010010010010,
        //tile_code 167
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000011011011011011011011011000000001,
        48'b000000000000011011011011011011011011011011011011,
        48'b000000000011100100100100100100100100100011011011,
        48'b010010010011100100100100100100100100100100100100,
        //tile_code 168
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b011011000000000000000001000000000000000000000001,
        48'b011011011011011011011011011011011000000000000001,
        48'b100011011011011011011011011011011011011011010010,
        //tile_code 169
        48'b000000000001001000000001001000000001001000000001,
        48'b001010010010011010010010011010010010011010010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        //tile_code 170
        48'b000001001000000001001000000001001000000001001000,
        48'b010011011011010011011011010011011011010011011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        //tile_code 171
        48'b000001001000000001001000000001001000000001001001,
        48'b010011011011010011011011010011011011010011011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        //tile_code 172
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        //tile_code 173
        48'b000001001001001001001001001001001001001001001000,
        48'b001010010001001000001001001001000001001010010001,
        48'b001010001000010001011011011011001000010001010001,
        48'b001001000010001011011011011011011001000010001001,
        48'b001000010000001011010010010010011001010000010001,
        48'b001000000010001010010010010010010001000010000001,
        48'b001000000000010001010010010010001000010000000001,
        48'b001001000011000010001001001001010000011000001001,
        48'b001000001000011000010000010000011000011001000001,
        48'b001011000001001000011000011000011001001000011001,
        48'b001011011000001001001001001001001001000011011001,
        48'b001011001001011011011011011011011011001001011001,
        48'b001001000000000000000000000000000000000000001001,
        48'b001011011011011011011011011011011011011011011001,
        48'b001011011011011011011011011011011011011011011001,
        48'b000001001001001001001001001001001001001001001000,
        //tile_code 174
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile_code 175
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        //tile_code 176
        48'b000001010011011001010011011001010011011001010011,
        48'b000001010011011001010011011001010011011001010011,
        48'b000000000011011000000011011000000011011000000011,
        48'b000011011000000011011000000011011000000011011000,
        48'b000001010011011001010011011001010011011001010011,
        48'b000001010011011001010011011001010011011001010011,
        48'b000000000011011000000011011000000011011000000011,
        48'b000011011000000011011000000011011000000011011000,
        48'b000001010011011001010011011001010011011001010011,
        48'b000001010011011001010011011001010011011001010011,
        48'b000000000011011000000011011000000011011000000011,
        48'b000011011000000011011000000011011000000011011000,
        48'b000001010011011001010011011001010011011001010011,
        48'b000001010011011001010011011001010011011001010011,
        48'b000000000011011000000011011000000011011000000011,
        48'b000011011000000011011000000011011000000011011000,
        //tile_code 177
        48'b000001010000000001010000000001010000000001010000,
        48'b000001010000000001010000000001010000000001010000,
        48'b000011011000000011011000000011011000000011011000,
        48'b011000000011011000000011011000000011011000000011,
        48'b000001010000000001010000000001010000000001010000,
        48'b000001010000000001010000000001010000000001010000,
        48'b000011011000000011011000000011011000000011011000,
        48'b011000000011011000000011011000000011011000000011,
        48'b000001010000000001010000000001010000000001010000,
        48'b000001010000000001010000000001010000000001010000,
        48'b000011011000000011011000000011011000000011011000,
        48'b011000000011011000000011011000000011011000000011,
        48'b000001010000000001010000000001010000000001010000,
        48'b000001010000000001010000000001010000000001010000,
        48'b000011011000000011011000000011011000000011011000,
        48'b011000000011011000000011011000000011011000000011,
        //tile_code 178
        48'b000001010000000001010000000001010000000001010011,
        48'b000001010000000001010000000001010000000001010011,
        48'b000011011000000011011000000011011000000011011011,
        48'b011000000011011000000011011000000011011000000011,
        48'b000001010000000001010000000001010000000001010011,
        48'b000001010000000001010000000001010000000001010011,
        48'b000011011000000011011000000011011000000011011011,
        48'b011000000011011000000011011000000011011000000011,
        48'b000001010000000001010000000001010000000001010011,
        48'b000001010000000001010000000001010000000001010011,
        48'b000011011000000011011000000011011000000011011011,
        48'b011000000011011000000011011000000011011000000011,
        48'b000001010000000001010000000001010000000001010011,
        48'b000001010000000001010000000001010000000001010011,
        48'b000011011000000011011000000011011000000011011011,
        48'b011000000011011000000011011000000011011000000011,
        //tile_code 179
        48'b000001001001001001001001001001001001001001001001,
        48'b001010010010010010010010010010010010010010010010,
        48'b001010011000000000000000000000000000000000000000,
        48'b001010000011011011011011011011011011011011011011,
        48'b001010000000000000000000000000000000000000000000,
        48'b001010000011011011011011011011011011011011011011,
        48'b001010000011011011011011011011011011011011011011,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        //tile_code 180
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        //tile_code 181
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010000,
        48'b001001001001001001001001001001001001001011010000,
        48'b011011011011011011011011011011011011011001010000,
        48'b001001001001001001001001001001001001001001010000,
        48'b011011011011011011011011011011011011011001010000,
        48'b011011011011011011011011011011011011011001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        //tile_code 182
        48'b000000001001001001001001001010010010010010010010,
        48'b000000001001001001001001001010010010010010010010,
        48'b000000001001001001001001001010001001010010011010,
        48'b000000001001001001001001001010010001001001001001,
        48'b000000001001001001001001001001010000000000001001,
        48'b000000001001001001001001001001010010000100100101,
        48'b000000001001001001001001001001010010011010100100,
        48'b000000001001001001001001001001001010010011010100,
        48'b000000001001001001001001001001001010010010011000,
        48'b000000001001001001001001001001001001010010010010,
        48'b000000001001001001001001001001001001010010010010,
        48'b000000001001001001001001001001001001001010010010,
        48'b000000001001001001001001001001001001001001010010,
        48'b000000001001001001001001001001001001001001001001,
        48'b000000001001001001001001001001001001001001001001,
        48'b000000001001001001001001001001001001001001001001,
        //tile_code 183
        48'b000000000000001001001001001001001000001001000000,
        48'b010000000000000000000000000000000000001000001001,
        48'b010010000000000000000000000000000000000001001001,
        48'b011010100000000000000000000000000000000000001001,
        48'b011010100000000000000000001001001000000000000000,
        48'b101010100000001101101000001000000000000000000001,
        48'b000100100000100100101101000000000000000000000000,
        48'b000000000000100100100000000000000000000000000000,
        48'b100000000000000000000000000000000100100100000000,
        48'b010010000000000000000000000100100100011000000000,
        48'b010010010100100100100100100010010010000000100100,
        48'b010010010010010010010010010010010010000000100101,
        48'b010010010010010010010010010010101101000000000101,
        48'b010010010010010010010010101101101101000000000000,
        48'b101101101101101101101101101101101100000000000000,
        48'b101101101101101101101101101101101000000000000000,
        //tile_code 184
        48'b000000000000000000000001001001000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001010010001001001001000001001001001001,
        48'b000001001001010010001001001000000000001001001001,
        48'b001000000000000000000011011011000000001001001001,
        48'b000000000000000010100100100100100000000001100011,
        48'b000000000000000010100100100100100100100010100100,
        48'b000001001000001010100100100100100100010010010100,
        48'b000001000001001010010100100100000000000000100100,
        48'b001000001001001001001100100100100000000000000000,
        48'b000001000001000001001001010100100000000010010000,
        48'b100100100000001000001001010000000000000010010000,
        48'b100100100100000000000000000000000000000000000000,
        48'b010100100100100010000000000000000000000000000000,
        48'b000000010100100010000000000000000000000000000011,
        48'b000000000000000000000000000000000000000000011011,
        //tile_code 185
        48'b000000000000000001010010010010010010010010010010,
        48'b000000000000000000010010010010010010010010010010,
        48'b000000000000000000000000010010010010010010010010,
        48'b000000000000000000000000000001000010010010010010,
        48'b000000000000000000000000000000001001001010010010,
        48'b011000000000000000000000000000000000001001001001,
        48'b100011010000000000000000000000000000000000000000,
        48'b100100000000000000000000000000010010010010010010,
        48'b100001000000000000000000010010010011011011011011,
        48'b001001001000000000000010010011011011011100100100,
        48'b001001000000000001001100100100100100100100100100,
        48'b001000001001001011011100100100100100100100100100,
        48'b001001000011100100100100100100100100100100100100,
        48'b001011100100100100100100100100100100100100100100,
        48'b011100100100100100100100100100100100100100100100,
        48'b100100100100100100100100100100100100100100100100,
        //tile_code 186
        48'b000000000000000001001001001001001010001001001001,
        48'b000000000000000000000001001001001010001001001001,
        48'b000000000000000000000000000001001011011011011011,
        48'b000000000000000000000011011011011011100011011011,
        48'b000000000000000011011011011011011011011011011011,
        48'b011011011011011011011011011000000011100100100000,
        48'b100100100100100100100100100000000100100011011101,
        48'b000100100100100100100100100100100011011101101101,
        48'b000000000000000000000000000000110110110101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        //tile_code 187
        48'b000000000001010010010010010010010010010010010010,
        48'b000000000010010010010010010010010010010010010010,
        48'b011011011011011010010010010010010010010010100100,
        48'b011011011011010010010101101101101101101101010010,
        48'b011010010010010101101101101101101101101101101101,
        48'b010010110110110110110110110110110110110110110110,
        48'b110110110110110110110110110110110110110110110110,
        48'b110110110110110110110110110110110110110110101101,
        48'b110110110110110110110110110110110110101101101101,
        48'b110110110110110110110110110110101101101101101101,
        48'b110110110110110110110110110101101101101101101101,
        48'b110110110110110110110110101101101101101101101010,
        48'b110110110110110110110110101101101101101101101010,
        48'b110110110110110110110110101101101101101101101101,
        48'b110110110110110110110110110110110110110110110110,
        48'b110110110110110110110110110110110110110110110110,
        //tile_code 188
        48'b000001001001001001010010010010010010001001001001,
        48'b000001001001001001010010010010010010010010010010,
        48'b001001001001001001010010010010010010010010010010,
        48'b000000000000000000000010010010010010010010010000,
        48'b011011011011011011011011010010010010010010010000,
        48'b100100100011011011011011011010001010010010010000,
        48'b011011011011011011010010010010001010010010010010,
        48'b011011011011011010010010010010010010010010010010,
        48'b011011011000000010010010010010010010010100100000,
        48'b011011011010010010010010010010010010010000100000,
        48'b011000010010010010010010010010010010010010010010,
        48'b000010010010010010010010010010010010010010010010,
        48'b000010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b100100100100100100100100100100100100100100100100,
        48'b100100100100100100100100100100100100100100100100,
        //tile_code 189
        48'b000001001001001001001001000000000000000000000000,
        48'b001001001001001001001001001000000000000000000000,
        48'b001001001001001001001001001001000000010000000000,
        48'b011011100100100001001001001001000000000000000000,
        48'b011011011011011010001001001000000000000000000000,
        48'b010010010010010001001001001000000000000000000001,
        48'b001001001001001001001001010001001001001010001010,
        48'b001001001001001001001001001001001001001010001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001010010010,
        48'b001001001001001001001001001001001001010100011100,
        48'b001001001001001001001001001001001010010100011011,
        48'b010010010010010010010010010010010010100100011011,
        48'b011011011011011011011011011011011011100100011011,
        48'b011011011011011011011011011011011011011011100011,
        //tile_code 190
        48'b000000001001001001001010010010010010010010010010,
        48'b000000010011001001001001001001011011011010010010,
        48'b000000010010011001001001001001001001011000000010,
        48'b000100000010010010010010001001001001000000000000,
        48'b100100100000000000000000000000000000000000000000,
        48'b100100100100000000000000000000000000000000000000,
        48'b100100100100000000000000000000000000000000000000,
        48'b100100100100000000000000000000000000100100100100,
        48'b100100100000100100100100100100100100100100100100,
        48'b100000000100010010010010010010010010010010010010,
        48'b010010010010010011011001001001001001001001001001,
        48'b011011011011011011011011001001001001001001001001,
        48'b001001001001001001001001011001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        //tile_code 191
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001000000,
        48'b001001001001001001001001001001001000000000010010,
        48'b011011011011011011011011011011000000100100010010,
        48'b011011011011011011011011011011000100010010010010,
        48'b000000000000000000000011011000000100010010010010,
        48'b010010010010010100000000000000100010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        //tile_code 192
        48'b000000001001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000001001001001001001001001001001001,
        48'b010010010010010000001001001001001001001001001001,
        48'b010010010010010010000001001001001001001001001001,
        48'b010010010010010010011000001001001001100100001001,
        48'b010010010010010010011000000000000000000100100100,
        48'b010010010010010010010011011011011010000000000100,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        //tile_code 193
        48'b000000000000000000000000000000001001001001001001,
        48'b000000000000000000000000000000000000001001000000,
        48'b000000000000000000000000000000000000000000000010,
        48'b000000000000000000000000000000000000000000000010,
        48'b000000000000000000000000000000000000000000000010,
        48'b000000000000000000000010010010010010010010010010,
        48'b000000000000000000010010010010010010010010010010,
        48'b000000000000000010010010010010010010010010010010,
        48'b000000000000010010010010000000000000000000010010,
        48'b010000000000010010010000000000000000000000000010,
        48'b010010010010010010000010000000000000000000010000,
        48'b001001010010010010010000010010000010000010000010,
        48'b011001001010010010010010010000010010010000010010,
        48'b100011001001001001001001010010010010010010010010,
        48'b100100011011011011001001001001001001010010010010,
        48'b100100100100100100011011011011011011001001001001,
        //tile_code 194
        48'b000000000000001010010010000000000011100100100100,
        48'b010000000001001001001001000000101000000000110110,
        48'b001001001001001110000000101101101101101101101101,
        48'b110110001001110110101101101101101101101101101101,
        48'b101110110001101101101101101101101101101101101101,
        48'b101101101101101101101101110101101101101000000101,
        48'b101101101101101101101101101101101000000000101000,
        48'b101101101101101101101101101101101000000000000101,
        48'b101101101101101101101101101101000000101000101101,
        48'b101101101101101101101101101000000101000101000101,
        48'b101101101101101101101110101101101000101000101101,
        48'b101101101101101101101101101101101101101101101110,
        48'b101101101101101101101101101101101101101101110110,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b110101101101101101101101101101101101101101101101,
        //tile_code 195
        48'b000000000001010010010010010010010011011011011011,
        48'b001001001010010010011011011011011011011011011011,
        48'b001001001010010010011011011011011011011011011011,
        48'b100101001010010010010011011011011011011011011011,
        48'b100100001010010010010011011011011011011011011011,
        48'b100100001010010010010010011011011011011011011011,
        48'b100100001010010010010010010011011011011011011011,
        48'b100100001001010010010010010011011011011011011011,
        48'b100100100001001010010010010010011011011011011011,
        48'b100100100100001001001010010010010011011011011011,
        48'b100100100100100001001001010010010010011011011011,
        48'b100100100100100100100001001010010010010011011011,
        48'b100100100100100100100001010010010010010010011011,
        48'b100100100100001001001010010011011011011011011011,
        48'b100100001001010010010010011011011011011011011011,
        48'b001001010010010010011011011011011011011011011011,
        //tile_code 196
        48'b000000000000000000000000000000000000001001001001,
        48'b000000000000000000000000000000000000001001001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        //tile_code 197
        48'b000001001001001001001001001001001001001001001001,
        48'b001010010010010010010010010010010010010010010010,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        //tile_code 198
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        //tile_code 199
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        //tile_code 200
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        //tile_code 201
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        //tile_code 202
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011
    };

    assign data = ROM[addr];

endmodule