module car_rom (
    input  logic [3:0] Tile,
    input  logic [5:0] PixelX,
    input  logic [4:0] PixelY,
    output logic [5:0] Data
);

    logic [51:0] data;
    logic [8:0] bitmapIdx;
    logic [143:0] bitmap;
    logic [2:0] color;

    localparam bit [51:0] DATA [16] = '{


        // <--- FILE: ASSETS\CAR\BLUE.PNG --->

        //tile 0
        52'b0001110100010100100100111000100010011101110000000000,
        //tile 1
        52'b0001110100010100100100111000100010011101110000000001,
        //tile 2
        52'b0001110100010100100100111000100010011101110000000010,
        //tile 3
        52'b0001110100010100100100111000100010011101110000000011,

        // <--- FILE: ASSETS\CAR\GREEN.PNG --->

        //tile 0
        52'b0001110010011000100101000110010101011110000000000100,
        //tile 1
        52'b0001110010011000100101000110010101011110000000000101,
        //tile 2
        52'b0001110010011000100101000110010101011110000000000110,
        //tile 3
        52'b0001110010011000100101000110010101011110000000000111,

        // <--- FILE: ASSETS\CAR\RED.PNG --->

        //tile 0
        52'b0001110010011000100111000111011110010110110000001000,
        //tile 1
        52'b0001110010011000100111000111011110010110110000001001,
        //tile 2
        52'b0001110010011000100111000111011110010110110000001010,
        //tile 3
        52'b0001110010011000100111000111011110010110110000001011,

        // <--- FILE: ASSETS\CAR\YELLOW.PNG --->

        //tile 0
        52'b0001111110110010011001010101101110101000100000001100,
        //tile 1
        52'b0001111110110010011001010101101110101000100000001101,
        //tile 2
        52'b0001111110110010011001010101101110101000100000001110,
        //tile 3
        52'b0001111110110010011001010101101110101000100000001111
    
    };

    localparam bit [143:0] BITMAPS [416] = '{


        // <--- FILE: ASSETS\CAR\BLUE.PNG --->

        //tile 0, VRAM 52'b0001110100010100100100111000100010011101110000000000
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000,
        144'b000000000000000000000000000000000000000000000000000000000001001010011011011011011011011011011011011011011011011011011011011011011011011011010000,
        144'b000000000000000000000000000000000000000000000000000000001100100011001001001001001001001001001001001001001001001001001001001001001001001001011001,
        144'b000000000000000000000000000000000000000000000000000001100100101101011011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b000000000000000000000000000000000000000000000000001100011100101011010010010010010010010010010010011101101101101101101101101101101101101101101001,
        144'b000001001001001001001001001001001001001001001001100011011100101011010011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100100100100100100100100100100100100100100100011010011100101011010011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100101001001001001001001001001001001001001110011010011100101011001011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100001110110110110110110110110110110110110110011011011100101011001011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100001100100100100100100100100100100100100110011011011100101011001011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100001100101101101101101101101101101101101110011011011100101011001001001001001001001001001001001001001001001001001001001001001001001001101001,
        144'b001100001100101101101101101101101101101101101110011011011100100001011011011011011011011011011011011011011011011011011011011011011011011011001001,
        144'b001100001100101101101101101101101101101101101110011011101001001011001001001001001001001001001001001001001001001001001001001001001001001001011001,
        144'b001100001100100100100101101101101101101101101110011101001100100100100100100100100100100100100100100100100100100100100100100100100100100100100001,
        144'b001100001001001001001001001001001001001001001110110001100001011001011011011011011011011011101011001011011011011011011011101011001011011011101001,
        144'b001100101101101101101101101101101101101101101110001101101001011001011011011011011011011011101011001011011011011011011011101011001011011011101001,
        144'b001001001001001001001001001001001001001001001001100001001001110110110110110110110110110110001110110110110110110110110110001101101101101101101001,
        144'b001100100100100100100100100100100100100100100100100101101001110100100100100100100011011100001110100100100100100011011100001101101101101101101001,
        144'b001101101101101101101101101101101101101101101101101101101001110100101101101101101101101101001110100101101101101101101101001101101101101101101001,
        144'b001101101101101101101001001001001001001001001001001101101001110100100100101101101101101101001001001001001001001001001001001101101101101101101001,
        144'b000001001001001001001001100101101101101101101110001001001001001001001001001001001001001001001001100101101101101101101110001001001001001001001001,
        144'b000001101101101101110011011011011011011011011011011110101101101101101101101101101101101101110011011011011011011011011011011110101101101101001000,
        144'b000000011011011011011111001111001111001111111111111011011011011011011011011011011011011011011111001111001111001111111111111011011011011011111000,
        144'b000000111111111111111011011001001001001001001011011111111111111111111111111111111111111111111011011001001001001001001011011111111111111111111000,
        144'b000000000111111111111111111011011011011011011111111111111111111111111111111111111111111111111111111011011011011011011111111111111111111111000000,
        //tile 1, VRAM 52'b0001110100010100100100111000100010011101110000000001
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000,
        144'b000000000000000000000000000000000000000000000000000000000001001010011011011011011011011011011011011011011011011011011011011011011011011011010000,
        144'b000000000000000000000000000000000000000000000000000000001100100011001001001001001001001001001001001001001001001001001001001001001001001001011001,
        144'b000000000000000000000000000000000000000000000000000001100100101101011011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b000000000000000000000000000000000000000000000000001100011100101011010010010010010010010010010010011101101101101101101101101101101101101101101001,
        144'b000001001001001001001001001001001001001001001001100011011100101011010011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100100100100100100100100100100100100100100100011010011100101011010011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100101001001001001001001001001001001001001110011010011100101011001011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100001110110110110110110110110110110110110110011011011100101011001011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100001100100100100100100100100100100100100110011011011100101011001011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100001100101101101101101101101101101101101110011011011100101011001001001001001001001001001001001001001001001001001001001001001001001001101001,
        144'b001100001100101101101101101101101101101101101110011011011100100001011011011011011011011011011011011011011011011011011011011011011011011011001001,
        144'b001100001100101101101101101101101101101101101110011011101001001011001001001001001001001001001001001001001001001001001001001001001001001001011001,
        144'b001100001100100100100101101101101101101101101110011101001100100100100100100100100100100100100100100100100100100100100100100100100100100100100001,
        144'b001100001001001001001001001001001001001001001110110001100001011001011011011011011011011011101011001011011011011011011011101011001011011011101001,
        144'b001100101101101101101101101101101101101101101110001101101001011001011011011011011011011011101011001011011011011011011011101011001011011011101001,
        144'b001001001001001001001001001001001001001001001001100001001001110110110110110110110110110110001110110110110110110110110110001101101101101101101001,
        144'b001100100100100100100100100100100100100100100100100101101001110100100100100100100011011100001110100100100100100011011100001101101101101101101001,
        144'b001101101101101101101101101101101101101101101101101101101001110100101101101101101101101101001110100101101101101101101101001101101101101101101001,
        144'b001101101101101101101001001001001001001001001001001101101001110100100100101101101101101101001001001001001001001001001001001101101101101101101001,
        144'b000001001001001001001001100101101101101101101110001001001001001001001001001001001001001001001001100101101101101101101110001001001001001001001001,
        144'b000001101101101101110011011011011011011011011011011110101101101101101101101101101101101101110011011011011011011011011011011110101101101101001000,
        144'b000000011011011011011111111111001111001111001111111011011011011011011011011011011011011011011111111111001111001111001111111011011011011011111000,
        144'b000000111111111111111011011001001001001001001011011111111111111111111111111111111111111111111011011001001001001001001011011111111111111111111000,
        144'b000000000111111111111111111011011011011011011111111111111111111111111111111111111111111111111111111011011011011011011111111111111111111111000000,
        //tile 2, VRAM 52'b0001110100010100100100111000100010011101110000000010
        144'b000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000,
        144'b000000000000000000000000000000000000000000000000000000000001001010011011011011011011011011011011011011011011011011011011011011011011011011010000,
        144'b000000000000000000000000000000000000000000000000000000001100100011001001001001001001001001001001001001001001001001001001001001001001001001011001,
        144'b000000000000000000000000000000000000000000000000000001100100101101011011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b000000000000000000000000000000000000000000000000001100011100101011010010010010010010010010010010011101101101101101101101101101101101101101101001,
        144'b000001001001001001001001001001001001001001001001100011011100101011010011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100100100100100100100100100100100100100100100011010011100101011010011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100101001001001001001001001001001001001001110011010011100101011001011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100001110110110110110110110110110110110110110011011011100101011001011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100001100100100100100100100100100100100100110011011011100101011001011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100001100101101101101101101101101101101101110011011011100101011001001001001001001001001001001001001001001001001001001001001001001001001101001,
        144'b001100001100101101101101101101101101101101101110011011011100100001011011011011011011011011011011011011011011011011011011011011011011011011001001,
        144'b001100001100101101101101101101101101101101101110011011101001001011001001001001001001001001001001001001001001001001001001001001001001001001011001,
        144'b001100001100100100100101101101101101101101101110011101001100100100100100100100100100100100100100100100100100100100100100100100100100100100100001,
        144'b001100001001001001001001001001001001001001001110110001100001011001011011011011011011011011101011001011011011011011011011101011001011011011101001,
        144'b001100101101101101101101101101101101101101101110001101101001011001011011011011011011011011101011001011011011011011011011101011001011011011101001,
        144'b001001001001001001001001001001001001001001001001100001001001110110110110110110110110110110001110110110110110110110110110001101101101101101101001,
        144'b001100100100100100100100100100100100100100100100100101101001110100100100100100100011011100001110100100100100100011011100001101101101101101101001,
        144'b001101101101101101101101101101101101101101101101101101101001110100101101101101101101101101001110100101101101101101101101001101101101101101101001,
        144'b001101101101101101101001001001001001001001001001001101101001110100100100101101101101101101001001001001001001001001001001001101101101101101101001,
        144'b000001001001001001001001100101101101101101101110001001001001001001001001001001001001001001001001100101101101101101101110001001001001001001001001,
        144'b000001101101101101110011011011011011011011011011011110101101101101101101101101101101101101110011011011011011011011011011011110101101101101001000,
        144'b000000011011011011011111001111001111001111111111111011011011011011011011011011011011011011011111001111001111001111111111111011011011011011111000,
        144'b000000111111111111111011011001001001001001001011011111111111111111111111111111111111111111111011011001001001001001001011011111111111111111111000,
        144'b000000111111111111111011011001001001001001001011011111111111111111111111111111111111111111111011011001001001001001001011011111111111111111111000,
        144'b000000000111111111111111111011011011011011011111111111111111111111111111111111111111111111111111111011011011011011011111111111111111111111000000,
        //tile 3, VRAM 52'b0001110100010100100100111000100010011101110000000011
        144'b000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000,
        144'b000000000000000000000000000000000000000000000000000000000001001010011011011011011011011011011011011011011011011011011011011011011011011011010000,
        144'b000000000000000000000000000000000000000000000000000000001100100011001001001001001001001001001001001001001001001001001001001001001001001001011001,
        144'b000000000000000000000000000000000000000000000000000001100100101101011011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b000000000000000000000000000000000000000000000000001100011100101011010010010010010010010010010010011101101101101101101101101101101101101101101001,
        144'b000001001001001001001001001001001001001001001001100011011100101011010011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100100100100100100100100100100100100100100100011010011100101011010011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100101001001001001001001001001001001001001110011010011100101011001011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100001110110110110110110110110110110110110110011011011100101011001011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100001100100100100100100100100100100100100110011011011100101011001011011011011011011011011011011101101101101101101101101101101101101101101001,
        144'b001100001100101101101101101101101101101101101110011011011100101011001001001001001001001001001001001001001001001001001001001001001001001001101001,
        144'b001100001100101101101101101101101101101101101110011011011100100001011011011011011011011011011011011011011011011011011011011011011011011011001001,
        144'b001100001100101101101101101101101101101101101110011011101001001011001001001001001001001001001001001001001001001001001001001001001001001001011001,
        144'b001100001100100100100101101101101101101101101110011101001100100100100100100100100100100100100100100100100100100100100100100100100100100100100001,
        144'b001100001001001001001001001001001001001001001110110001100001011001011011011011011011011011101011001011011011011011011011101011001011011011101001,
        144'b001100101101101101101101101101101101101101101110001101101001011001011011011011011011011011101011001011011011011011011011101011001011011011101001,
        144'b001001001001001001001001001001001001001001001001100001001001110110110110110110110110110110001110110110110110110110110110001101101101101101101001,
        144'b001100100100100100100100100100100100100100100100100101101001110100100100100100100011011100001110100100100100100011011100001101101101101101101001,
        144'b001101101101101101101101101101101101101101101101101101101001110100101101101101101101101101001110100101101101101101101101001101101101101101101001,
        144'b001101101101101101101001001001001001001001001001001101101001110100100100101101101101101101001001001001001001001001001001001101101101101101101001,
        144'b000001001001001001001001100101101101101101101110001001001001001001001001001001001001001001001001100101101101101101101110001001001001001001001001,
        144'b000001101101101101110011011011011011011011011011011110101101101101101101101101101101101101110011011011011011011011011011011110101101101101001000,
        144'b000000011011011011011111111111001111001111001111111011011011011011011011011011011011011011011111111111001111001111001111111011011011011011111000,
        144'b000000111111111111111011011001001001001001001011011111111111111111111111111111111111111111111011011001001001001001001011011111111111111111111000,
        144'b000000111111111111111011011001001001001001001011011111111111111111111111111111111111111111111011011001001001001001001011011111111111111111111000,
        144'b000000000111111111111111111011011011011011011111111111111111111111111111111111111111111111111111111011011011011011011111111111111111111111000000,

        // <--- FILE: ASSETS\CAR\GREEN.PNG --->

        //tile 4, VRAM 52'b0001110010011000100101000110010101011110000000000100
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000,
        144'b000000000000000000000000000000000000000001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001000000,
        144'b000000000000000000000000000000000000001010010011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011010001000,
        144'b000000000000000000000000000000000001010101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101010001,
        144'b000000001001001001001001001001001010101110101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101001,
        144'b000001010010010010010010010010010101110110101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101110101,
        144'b001010100001001001001001001001011101110101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101110101,
        144'b001010001011011011011011011011011101101101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010010010010010010010011101101101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010100100100100100100011101101101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010100100100100100100011101101101101011010010010010010100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010100100100100100100011101101100100001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001100101101,
        144'b001010001010010010100100100100011101100001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001100101,
        144'b001010100001001001001001001001011100001010010101101110101101110101101101101101101110101101101101110110101110101101101101101101101101100010001001,
        144'b001010100100100100100100100100011001101100100101110101101110110110101101101101110101101101110101101101110101101101101101110101110110101100010001,
        144'b001100001001001001001001001001001010011101101011011011011011011011011011011011011011011011011011011011011011011011011011011001011011011001001001,
        144'b001001110001010010010010010010010100011010010010010010010101101010011010010010010010101101010011010010010010010101101100100001100100100001110001,
        144'b001001001100010010010010010100100100011010100100100100100100100100011100100100100100100100100011100100100100100100100010011010010010010100001001,
        144'b001100100101101101101101101010010100011010010010100100100100100011010011010010010010010010011010011010010010010010010101101101101101101010100001,
        144'b001101101111111111111111111101101011001001001001001001001001001001001001001001001001001001001001001001001001001101101111111111111111111101101001,
        144'b101111111111110111110111110111111101011011011011011011011011011011011011011011011011011011011011011011011011011111111111110111110111110111111101,
        144'b101110110110111110111110111110110101101101101101101101101101101101101101101101101101101101101101101101101101101110110110111110111110111110110101,
        144'b000101101110110110110110110101101111111111111111111111111111111111111111111111111111111111111111111111111111111101101110110110110110110101101000,
        144'b000111111101101101101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101101101101101111111000,
        //tile 5, VRAM 52'b0001110010011000100101000110010101011110000000000101
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000,
        144'b000000000000000000000000000000000000000001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001000000,
        144'b000000000000000000000000000000000000001010010011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011010001000,
        144'b000000000000000000000000000000000001010101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101010001,
        144'b000000001001001001001001001001001010101110101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101001,
        144'b000001010010010010010010010010010101110110101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101110101,
        144'b001010100001001001001001001001011101110101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101110101,
        144'b001010001011011011011011011011011101101101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010010010010010010010011101101101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010100100100100100100011101101101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010100100100100100100011101101101101011010010010010010100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010100100100100100100011101101100100001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001100101101,
        144'b001010001010010010100100100100011101100001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001100101,
        144'b001010100001001001001001001001011100001010010101101110101101110101101101101101101110101101101101110110101110101101101101101101101101100010001001,
        144'b001010100100100100100100100100011001101100100101110101101110110110101101101101110101101101110101101101110101101101101101110101110110101100010001,
        144'b001100001001001001001001001001001010011101101011011011011011011011011011011011011011011011011011011011011011011011011011011001011011011001001001,
        144'b001001110001010010010010010010010100011010010010010010010101101010011010010010010010101101010011010010010010010101101100100001100100100001110001,
        144'b001001001100010010010010010100100100011010100100100100100100100100011100100100100100100100100011100100100100100100100010011010010010010100001001,
        144'b001100100101101101101101101010010100011010010010100100100100100011010011010010010010010010011010011010010010010010010101101101101101101010100001,
        144'b001101101111111111111111111101101011001001001001001001001001001001001001001001001001001001001001001001001001001101101111111111111111111101101001,
        144'b101111111111110111110111111111111101011011011011011011011011011011011011011011011011011011011011011011011011011111111111110111110111111111111101,
        144'b101111111110111110111110110110110101101101101101101101101101101101101101101101101101101101101101101101101101101111111110111110111110110110110101,
        144'b000101101111110110110110110101101111111111111111111111111111111111111111111111111111111111111111111111111111111101101111110110110110110101101000,
        144'b000111111101101101101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101101101101101111111000,
        //tile 6, VRAM 52'b0001110010011000100101000110010101011110000000000110
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000,
        144'b000000000000000000000000000000000000000001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001000000,
        144'b000000000000000000000000000000000000001010010011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011010001000,
        144'b000000000000000000000000000000000001010101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101010001,
        144'b000000001001001001001001001001001010101110101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101001,
        144'b000001010010010010010010010010010101110110101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101110101,
        144'b001010100001001001001001001001011101110101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101110101,
        144'b001010001011011011011011011011011101101101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010010010010010010010011101101101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010100100100100100100011101101101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010100100100100100100011101101101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010100100100100100100011101101100100001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001100101101,
        144'b001010001010010010100100100100011101100001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001100101,
        144'b001010100001001001001001001001011100001010010101101110101101110101101101101101101110101101101101110110101110101101101101101101101101100010001001,
        144'b001010100100100100100100100100011001101100100101110101101110110110101101101101110101101101110101101101110101101101101101110101110110101100010001,
        144'b001100001001001001001001001001001010011101101011011011011011011011011011011011011011011011011011011011011011011011011011011001011011011001001001,
        144'b001001110001010010010010010010010100011010010010010010010101101010011010010010010010101101010011010010010010010101101100100001100100100001110001,
        144'b001001001100010010010010010100100100011010100100100100100100100100011100100100100100100100100011100100100100100100100010011010010010010100001001,
        144'b001100100101101101101101101010010100011010010010100100100100100011010011010010010010010010011010011010010010010010010101101101101101101010100001,
        144'b001101101111111111111111111101101011001001001001001001001001001001001001001001001001001001001001001001001001001101101111111111111111111101101001,
        144'b101111111111110111110111111111111101011011011011011011011011011011011011011011011011011011011011011011011011011111111111110111110111111111111101,
        144'b101111111110111110111110110110110101101101101101101101101101101101101101101101101101101101101101101101101101101111111110111110111110110110110101,
        144'b000101101111110110110110110101101111111111111111111111111111111111111111111111111111111111111111111111111111111101101111110110110110110101101000,
        144'b000101101110111110111110111101101111111111111111111111111111111111111111111111111111111111111111111111111111111101101110111110111110111101101000,
        144'b000111111101101101101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101101101101101111111000,
        //tile 7, VRAM 52'b0001110010011000100101000110010101011110000000000111
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000,
        144'b000000000000000000000000000000000000000001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001000000,
        144'b000000000000000000000000000000000000001010010011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011010001000,
        144'b000000000000000000000000000000000001010101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101010001,
        144'b000000001001001001001001001001001010101110101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101001,
        144'b000001010010010010010010010010010101110110101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101110101,
        144'b001010100001001001001001001001011101110101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101110101,
        144'b001010001011011011011011011011011101101101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010010010010010010010011101101101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010100100100100100100011101101101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010100100100100100100011101101101101011010100100100100100100100100100100100100100100100100100100100100100100100100100100100011101101101,
        144'b001010001010100100100100100100011101101100100001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001100101101,
        144'b001010001010010010100100100100011101100001001010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010001100101,
        144'b001010100001001001001001001001011100001010010101101110101101110101101101101101101110101101101101110110101110101101101101101101101101100010001001,
        144'b001010100100100100100100100100011001101100100101110101101110110110101101101101110101101101110101101101110101101101101101110101110110101100010001,
        144'b001100001001001001001001001001001010011101101011011011011011011011011011011011011011011011011011011011011011011011011011011001011011011001001001,
        144'b001001110001010010010010010010010100011010010010010010010101101010011010010010010010101101010011010010010010010101101100100001100100100001110001,
        144'b001001001100010010010010010100100100011010100100100100100100100100011100100100100100100100100011100100100100100100100010011010010010010100001001,
        144'b001100100101101101101101101010010100011010010010100100100100100011010011010010010010010010011010011010010010010010010101101101101101101010100001,
        144'b001101101111111111111111111101101011001001001001001001001001001001001001001001001001001001001001001001001001001101101111111111111111111101101001,
        144'b101111111111110111110111110111111101011011011011011011011011011011011011011011011011011011011011011011011011011111111111110111110111110111111101,
        144'b101110110110110110111110111110110101101101101101101101101101101101101101101101101101101101101101101101101101101110110110110110111110111110110101,
        144'b000101101110110110110111110101101111111111111111111111111111111111111111111111111111111111111111111111111111111101101110110110110111110101101000,
        144'b000101101110110110111110111101101111111111111111111111111111111111111111111111111111111111111111111111111111111101101110110110111110111101101000,
        144'b000111111101101101101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101101101101101111111000,

        // <--- FILE: ASSETS\CAR\RED.PNG --->

        //tile 8, VRAM 52'b0001110010011000100111000111011110010110110000001000
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000001001010010010010010010010010010010010010010010010010001000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000001001010010011010100100100100100100100100100100100100100011010001000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000001001010010101101011010100100100100100100100100100100100100100011101010001001000000000000000,
        144'b000000000000001001001001001001001001001001001001001010010101101110101011010100100100100100100100100100100100100100011101101010010001001001001000,
        144'b000000001001010010010010010010010010010010010010010101101110110110101011010100100100100100100100100100100100100100011101110101101010010001010001,
        144'b000001010010001001001001001001001001001001001001011101110110110101101011010100100100100100100100100100100100100100011101110110110101011001010001,
        144'b001010100001011011011011011011011011011011011011011101110101101101101011010100100100100100100100100100100100100100011101101110110101011001010001,
        144'b001010001011010010010010010010010010010010010010011101101101101101101011010100100100100100100100100100100100100100011101101101101101011001010001,
        144'b001010001010100100100100100100100100100100100100011101101101101101101011010100100100100100100100100100100100100100011101101101101101011001010001,
        144'b001010001010100100100100100100100100100100100100011101101101101101101011010010010010010100100100100100100100100100011101101101101101011001010001,
        144'b001010001010100100100100100100100100100100100100011101101101101100100001001001001001001001001001001001001001001001001100101101101101011001010001,
        144'b001010001010010010010100100100100100100100100100011101101100100001001010010010010010010010010010010010010010010010010001100101101101011001010001,
        144'b001010001010001001001001001001001001001001001001011100100001001010010101101110101101110110110101101101101101101101101010001100100101011001010001,
        144'b001010001001100100100100100100100100100100100100011001001010101100100101110101101110110110101101101101101101101101101101010001001100011001010001,
        144'b001010100100001001001001001001001001001001001001001010010001011101101011011011011011011011001100100100100100100100100100001010010001001001001001,
        144'b001010001001010010010010010010010010010010010010010100100001011010010010010010010101101010001100100100100100100101101100001100100100001110011001,
        144'b001001110001100100100100100010010010010010010100100100100001011010100100100100100100100100001100100010010010010010010100001100100100100001001001,
        144'b001011001100100100100010010101101101101101101010010100100001011010010010100100100100100100001010010101101101101101101010001100011011100100100101,
        144'b000101011101011011011101101111111111111111111101101011011001001001001001001001001001001001011101101111111111111111111101101011011011011011011101,
        144'b000101011101011011101111111111110111110111110111111101011011011011011011011011011011011011101111111111110111110111110111111101011011011011101000,
        144'b000000101101101101101110110110111110111110111110110101101101101101101101101101101101101101101110110110111110111110111110110101101101101101111000,
        144'b000000111111111111111101101110110110110110110101101111111111111111111111111111111111111111111101101110110110110110110101101111111111111111111000,
        144'b000000000111111111111111111101101101101101101111111111111111111111111111111111111111111111111111111101101101101101101111111111111111111111000000,
        //tile 9, VRAM 52'b0001110010011000100111000111011110010110110000001001
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000001001010010010010010010010010010010010010010010010010001000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000001001010010011010100100100100100100100100100100100100100011010001000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000001001010010101101011010100100100100100100100100100100100100100011101010001001000000000000000,
        144'b000000000000001001001001001001001001001001001001001010010101101110101011010100100100100100100100100100100100100100011101101010010001001001001000,
        144'b000000001001010010010010010010010010010010010010010101101110110110101011010100100100100100100100100100100100100100011101110101101010010001010001,
        144'b000001010010001001001001001001001001001001001001011101110110110101101011010100100100100100100100100100100100100100011101110110110101011001010001,
        144'b001010100001011011011011011011011011011011011011011101110101101101101011010100100100100100100100100100100100100100011101101110110101011001010001,
        144'b001010001011010010010010010010010010010010010010011101101101101101101011010100100100100100100100100100100100100100011101101101101101011001010001,
        144'b001010001010100100100100100100100100100100100100011101101101101101101011010100100100100100100100100100100100100100011101101101101101011001010001,
        144'b001010001010100100100100100100100100100100100100011101101101101101101011010010010010010100100100100100100100100100011101101101101101011001010001,
        144'b001010001010100100100100100100100100100100100100011101101101101100100001001001001001001001001001001001001001001001001100101101101101011001010001,
        144'b001010001010010010010100100100100100100100100100011101101100100001001010010010010010010010010010010010010010010010010001100101101101011001010001,
        144'b001010001010001001001001001001001001001001001001011100100001001010010101101110101101110110110101101101101101101101101010001100100101011001010001,
        144'b001010001001100100100100100100100100100100100100011001001010101100100101110101101110110110101101101101101101101101101101010001001100011001010001,
        144'b001010100100001001001001001001001001001001001001001010010001011101101011011011011011011011001100100100100100100100100100001010010001001001001001,
        144'b001010001001010010010010010010010010010010010010010100100001011010010010010010010101101010001100100100100100100101101100001100100100001110011001,
        144'b001001110001100100100100100010010010010010010100100100100001011010100100100100100100100100001100100010010010010010010100001100100100100001001001,
        144'b001011001100100100100010010101101101101101101010010100100001011010010010100100100100100100001010010101101101101101101010001100011011100100100101,
        144'b000101011101011011011101101111111111111111111101101011011001001001001001001001001001001001011101101111111111111111111101101011011011011011011101,
        144'b000101011101011011101111111111110111110111111111111101011011011011011011011011011011011011101111111111110111110111111111111101011011011011101000,
        144'b000000101101101101101110110110111110111110110110110101101101101101101101101101101101101101101110110110111110111110110110110101101101101101111000,
        144'b000000111111111111111101101110110110110110110101101111111111111111111111111111111111111111111101101110110110110110110101101111111111111111111000,
        144'b000000000111111111111111111101101101101101101111111111111111111111111111111111111111111111111111111101101101101101101111111111111111111111000000,
        //tile 10, VRAM 52'b0001110010011000100111000111011110010110110000001010
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000001001010010010010010010010010010010010010010010010010001000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000001001010010011010100100100100100100100100100100100100100011010001000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000001001010010101101011010100100100100100100100100100100100100100011101010001001000000000000000,
        144'b000000000000001001001001001001001001001001001001001010010101101110101011010100100100100100100100100100100100100100011101101010010001001001001000,
        144'b000000001001010010010010010010010010010010010010010101101110110110101011010100100100100100100100100100100100100100011101110101101010010001010001,
        144'b000001010010001001001001001001001001001001001001011101110110110101101011010100100100100100100100100100100100100100011101110110110101011001010001,
        144'b001010100001011011011011011011011011011011011011011101110101101101101011010100100100100100100100100100100100100100011101101110110101011001010001,
        144'b001010001011010010010010010010010010010010010010011101101101101101101011010100100100100100100100100100100100100100011101101101101101011001010001,
        144'b001010001010100100100100100100100100100100100100011101101101101101101011010100100100100100100100100100100100100100011101101101101101011001010001,
        144'b001010001010100100100100100100100100100100100100011101101101101101101011010100100100100100100100100100100100100100011101101101101101011001010001,
        144'b001010001010100100100100100100100100100100100100011101101101101100100001001001001001001001001001001001001001001001001100101101101101011001010001,
        144'b001010001010010010010100100100100100100100100100011101101100100001001010010010010010010010010010010010010010010010010001100101101101011001010001,
        144'b001010001010001001001001001001001001001001001001011100100001001010010101101110101101110110110101101101101101101101101010001100100101011001010001,
        144'b001010001001100100100100100100100100100100100100011001001010101100100101110101101110110110101101101101101101101101101101010001001100011001010001,
        144'b001010100100001001001001001001001001001001001001001010010001011101101011011011011011011011001100100100100100100100100100001010010001001001001001,
        144'b001010001001010010010010010010010010010010010010010100100001011010010010010010010101101010001100100100100100100101101100001100100100001110011001,
        144'b001001110001100100100100100010010010010010010100100100100001011010100100100100100100100100001100100010010010010010010100001100100100100001001001,
        144'b001011001100100100100010010101101101101101101010010100100001011010010010100100100100100100001010010101101101101101101010001100011011100100100101,
        144'b000101011101011011011101101111111111111111111101101011011001001001001001001001001001001001011101101111111111111111111101101011011011011011011101,
        144'b000101011101011011101111111111110111110111111111111101011011011011011011011011011011011011101111111111110111110111111111111101011011011011101000,
        144'b000000101101101101101111111110111110110110111111111101101101101101101101101101101101101101101111111110111110110110111111111101101101101101111000,
        144'b000000111111111111111101101111110110110110110101101111111111111111111111111111111111111111111101101111110110110110110101101111111111111111111000,
        144'b000000111111111111111101101110111110110110110101101111111111111111111111111111111111111111111101101110111110110110110101101111111111111111111000,
        144'b000000000111111111111111111101101101101101101111111111111111111111111111111111111111111111111111111101101101101101101111111111111111111111000000,
        //tile 11, VRAM 52'b0001110010011000100111000111011110010110110000001011
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000001001010010010010010010010010010010010010010010010010001000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000001001010010011010100100100100100100100100100100100100100011010001000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000001001010010101101011010100100100100100100100100100100100100100011101010001001000000000000000,
        144'b000000000000001001001001001001001001001001001001001010010101101110101011010100100100100100100100100100100100100100011101101010010001001001001000,
        144'b000000001001010010010010010010010010010010010010010101101110110110101011010100100100100100100100100100100100100100011101110101101010010001010001,
        144'b000001010010001001001001001001001001001001001001011101110110110101101011010100100100100100100100100100100100100100011101110110110101011001010001,
        144'b001010100001011011011011011011011011011011011011011101110101101101101011010100100100100100100100100100100100100100011101101110110101011001010001,
        144'b001010001011010010010010010010010010010010010010011101101101101101101011010100100100100100100100100100100100100100011101101101101101011001010001,
        144'b001010001010100100100100100100100100100100100100011101101101101101101011010100100100100100100100100100100100100100011101101101101101011001010001,
        144'b001010001010100100100100100100100100100100100100011101101101101101101011010100100100100100100100100100100100100100011101101101101101011001010001,
        144'b001010001010100100100100100100100100100100100100011101101101101100100001001001001001001001001001001001001001001001001100101101101101011001010001,
        144'b001010001010010010010100100100100100100100100100011101101100100001001010010010010010010010010010010010010010010010010001100101101101011001010001,
        144'b001010001010001001001001001001001001001001001001011100100001001010010101101110101101110110110101101101101101101101101010001100100101011001010001,
        144'b001010001001100100100100100100100100100100100100011001001010101100100101110101101110110110101101101101101101101101101101010001001100011001010001,
        144'b001010100100001001001001001001001001001001001001001010010001011101101011011011011011011011001100100100100100100100100100001010010001001001001001,
        144'b001010001001010010010010010010010010010010010010010100100001011010010010010010010101101010001100100100100100100101101100001100100100001110011001,
        144'b001001110001100100100100100010010010010010010100100100100001011010100100100100100100100100001100100010010010010010010100001100100100100001001001,
        144'b001011001100100100100010010101101101101101101010010100100001011010010010100100100100100100001010010101101101101101101010001100011011100100100101,
        144'b000101011101011011011101101111111111111111111101101011011001001001001001001001001001001001011101101111111111111111111101101011011011011011011101,
        144'b000101011101011011101111111111110110110110111111111101011011011011011011011011011011011011101111111111110110110110111111111101011011011011101000,
        144'b000000101101101101101111111110111110110110110111111101101101101101101101101101101101101101101111111110111110110110110111111101101101101101111000,
        144'b000000111111111111111101101111110110110111110101101111111111111111111111111111111111111111111101101111110110110111110101101111111111111111111000,
        144'b000000111111111111111101101110111110111110111101101111111111111111111111111111111111111111111101101110111110111110111101101111111111111111111000,
        144'b000000000111111111111111111101101101101101101111111111111111111111111111111111111111111111111111111101101101101101101111111111111111111111000000,

        // <--- FILE: ASSETS\CAR\YELLOW.PNG --->

        //tile 12, VRAM 52'b0001111110110010011001010101101110101000100000001100
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000001010010010010010010010010010010001000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000001010001010010011011011011011011011001000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000001010001010010011011011011011011011001000000000000000000000000000000000000000000000000000000000,
        144'b000001001001001001001001001001001001001001001001010001001010010011011011011011011011001001001001001001001001001001001001001001001001001001000000,
        144'b001100100010010010010010010010010010010010010100001101001010010011011011011011011011001100100100100100100100100100100100100100100001001100001001,
        144'b001100100001001001001001001001001001001001001100001101001010010011011011011011011011001010010010010010010010010010010010010010010011001001001001,
        144'b001100001100100100100100100100100100100100100100001101001010010011011011011011011011001010010010010010010010010010010010010010010011001001001001,
        144'b001100001100100100100100100100100100100100100100001001001010010011011011011011011011001001001001001001001001001001001001001001001011001001001001,
        144'b001100001100100100100100100100100100100100100100001001001010010011011011011011011011001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100001001001010010010010011011011011011001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100001001100001001001001001001001001001001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100001100010001010010010010010010010010001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100100010001001010001001001001001001001001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100100100100011011011011011011011011100010001001001010001001001001001001001001100100100100011011011011011011011011011011011001001001001,
        144'b001001001001001001001001001001001001001001001001001001001001010001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        144'b001100100100100100100100100100100100100100100100100011001010010100100100100100010100001011011011011011011001001001001001001001001001101011001001,
        144'b001011011011011011011011011011011011011011011011011011001010010100011011011011011011001011011011011011011011011011011011011011011011001001011001,
        144'b001011011011011011011001001001001001001001001001001011001010010100100100011011011011001011011001001001001001001001001001001011011011011011011001,
        144'b001001001001001001001001100011011011011011011010001001001001001001001001001001001001001001001001100011011011011011011010001001001001001001001001,
        144'b000001011011011011010001001001001001001001001001001010011011011011011011011011011011011011010001001001001001001001001001001010011011011011001000,
        144'b000000001001001001001101101101111101111101111101101001001001001001001001001001001001001001001101101101111101111101111101101001001001001001111000,
        144'b000000111111111111111001001101101101101101101001001111111111111111111111111111111111111111111001001101101101101101101001001111111111111111111000,
        144'b000000000111111111111111111001001001001001001111111111111111111111111111111111111111111111111111111001001001001001001111111111111111111111000000,
        //tile 13, VRAM 52'b0001111110110010011001010101101110101000100000001101
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000001010010010010010010010010010010001000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000001010001010010011011011011011011011001000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000001010001010010011011011011011011011001000000000000000000000000000000000000000000000000000000000,
        144'b000001001001001001001001001001001001001001001001010001001010010011011011011011011011001001001001001001001001001001001001001001001001001001000000,
        144'b001100100010010010010010010010010010010010010100001101001010010011011011011011011011001100100100100100100100100100100100100100100001001100001001,
        144'b001100100001001001001001001001001001001001001100001101001010010011011011011011011011001010010010010010010010010010010010010010010011001001001001,
        144'b001100001100100100100100100100100100100100100100001101001010010011011011011011011011001010010010010010010010010010010010010010010011001001001001,
        144'b001100001100100100100100100100100100100100100100001001001010010011011011011011011011001001001001001001001001001001001001001001001011001001001001,
        144'b001100001100100100100100100100100100100100100100001001001010010011011011011011011011001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100001001001010010010010011011011011011001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100001001100001001001001001001001001001001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100001100010001010010010010010010010010001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100100010001001010001001001001001001001001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100100100100011011011011011011011011100010001001001010001001001001001001001001100100100100011011011011011011011011011011011001001001001,
        144'b001001001001001001001001001001001001001001001001001001001001010001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        144'b001100100100100100100100100100100100100100100100100011001010010100100100100100010100001011011011011011011001001001001001001001001001101011001001,
        144'b001011011011011011011011011011011011011011011011011011001010010100011011011011011011001011011011011011011011011011011011011011011011001001011001,
        144'b001011011011011011011001001001001001001001001001001011001010010100100100011011011011001011011001001001001001001001001001001011011011011011011001,
        144'b001001001001001001001001100011011011011011011010001001001001001001001001001001001001001001001001100011011011011011011010001001001001001001001001,
        144'b000001011011011011010001001001001001001001001001001010011011011011011011011011011011011011010001001001001001001001001001001010011011011011001000,
        144'b000000001001001001001101101101111101111101101101101001001001001001001001001001001001001001001101101101111101111101101101101001001001001001111000,
        144'b000000111111111111111001001101101101101101101001001111111111111111111111111111111111111111111001001101101101101101101001001111111111111111111000,
        144'b000000000111111111111111111001001001001001001111111111111111111111111111111111111111111111111111111001001001001001001111111111111111111111000000,
        //tile 14, VRAM 52'b0001111110110010011001010101101110101000100000001110
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000001010010010010010010010010010010001000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000001010001010010011011011011011011011001000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000001010001010010011011011011011011011001000000000000000000000000000000000000000000000000000000000,
        144'b000001001001001001001001001001001001001001001001010001001010010011011011011011011011001001001001001001001001001001001001001001001001001001000000,
        144'b001100100010010010010010010010010010010010010100001101001010010011011011011011011011001100100100100100100100100100100100100100100001001100001001,
        144'b001100100001001001001001001001001001001001001100001101001010010011011011011011011011001010010010010010010010010010010010010010010011001001001001,
        144'b001100001100100100100100100100100100100100100100001101001010010011011011011011011011001010010010010010010010010010010010010010010011001001001001,
        144'b001100001100100100100100100100100100100100100100001001001010010011011011011011011011001001001001001001001001001001001001001001001011001001001001,
        144'b001100001100100100100100100100100100100100100100001001001010010011011011011011011011001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100001001001010010011011011011011011011001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100001001100001001001001001001001001001001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100001100010001010010010010010010010010001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100100010001001010001001001001001001001001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100100100100011011011011011011011011100010001001001010001001001001001001001001100100100100011011011011011011011011011011011001001001001,
        144'b001001001001001001001001001001001001001001001001001001001001010001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        144'b001100100100100100100100100100100100100100100100100011001010010100100100100100010100001011011011011011011001001001001001001001001001101011001001,
        144'b001011011011011011011011011011011011011011011011011011001010010100011011011011011011001011011011011011011011011011011011011011011011001001011001,
        144'b001011011011011011011001001001001001001001001001001011001010010100100100011011011011001011011001001001001001001001001001001011011011011011011001,
        144'b001001001001001001001001100011011011011011011010001001001001001001001001001001001001001001001001100011011011011011011010001001001001001001001001,
        144'b000001011011011011010001001001001001001001001001001010011011011011011011011011011011011011010001001001001001001001001001001010011011011011001000,
        144'b000000001001001001001111111101111101101101111111111001001001001001001001001001001001001001001111111101111101101101111111111001001001001001111000,
        144'b000000111111111111111001001111101101101101101001001111111111111111111111111111111111111111111001001111101101101101101001001111111111111111111000,
        144'b000000111111111111111001001101111101101101101001001111111111111111111111111111111111111111111001001101111101101101101001001111111111111111111000,
        144'b000000000111111111111111111001001001001001001111111111111111111111111111111111111111111111111111111001001001001001001111111111111111111111000000,
        //tile 15, VRAM 52'b0001111110110010011001010101101110101000100000001111
        144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000000001010010010010010010010010010010001000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000001010001010010011011011011011011011001000000000000000000000000000000000000000000000000000000000,
        144'b000000000000000000000000000000000000000000000000001010001010010011011011011011011011001000000000000000000000000000000000000000000000000000000000,
        144'b000001001001001001001001001001001001001001001001010001001010010011011011011011011011001001001001001001001001001001001001001001001001001001000000,
        144'b001100100010010010010010010010010010010010010100001101001010010011011011011011011011001100100100100100100100100100100100100100100001001100001001,
        144'b001100100001001001001001001001001001001001001100001101001010010011011011011011011011001010010010010010010010010010010010010010010011001001001001,
        144'b001100001100100100100100100100100100100100100100001101001010010011011011011011011011001010010010010010010010010010010010010010010011001001001001,
        144'b001100001100100100100100100100100100100100100100001001001010010011011011011011011011001001001001001001001001001001001001001001001011001001001001,
        144'b001100001100100100100100100100100100100100100100001001001010010011011011011011011011001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100001001001010010011011011011011011011001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100001001100001001001001001001001001001001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100001100010001010010010010010010010010001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100011011011011011011011011011011011100100010001001010001001001001001001001001110110110110110110110110110110110110110110011001001001001,
        144'b001011001100100100100011011011011011011011011100010001001001010001001001001001001001001100100100100011011011011011011011011011011011001001001001,
        144'b001001001001001001001001001001001001001001001001001001001001010001001001001001001001001001001001001001001001001001001001001001001001001001001001,
        144'b001100100100100100100100100100100100100100100100100011001010010100100100100100010100001011011011011011011001001001001001001001001001101011001001,
        144'b001011011011011011011011011011011011011011011011011011001010010100011011011011011011001011011011011011011011011011011011011011011011001001011001,
        144'b001011011011011011011001001001001001001001001001001011001010010100100100011011011011001011011001001001001001001001001001001011011011011011011001,
        144'b001001001001001001001001100011011011011011011010001001001001001001001001001001001001001001001001100011011011011011011010001001001001001001001001,
        144'b000001011011011011010001001001001001001001001001001010011011011011011011011011011011011011010001001001001001001001001001001010011011011011001000,
        144'b000000001001001001001111111101111101101101101111111001001001001001001001001001001001001001001111111101111101101101101111111001001001001001111000,
        144'b000000111111111111111001001111101101101111101001001111111111111111111111111111111111111111111001001111101101101111101001001111111111111111111000,
        144'b000000111111111111111001001101111101111101111001001111111111111111111111111111111111111111111001001101111101111101111001001111111111111111111000,
        144'b000000000111111111111111111001001001001001001111111111111111111111111111111111111111111111111111111001001001001001001111111111111111111111000000
    
    };

    always_comb
    begin
        data      = DATA[Tile];
        bitmapIdx = 9'd26 * data[3:0] + PixelY;
        bitmap    = BITMAPS[bitmapIdx];
        color     = bitmap[3*(47-PixelX) +: 3];
        Data      = data[6*color+4 +: 6];
    end

endmodule
