module text_rematch_rom (
    input  logic [8:0] PixelX,
    input  logic [5:0] PixelY,
    output logic [5:0] Data
);

    logic [47:0] data = 48'b00000000000000000000000000000111110101010000000;
    logic [5:0] bitmapIdx;
    logic [1196:0] bitmap;
    logic [2:0] color;

    localparam bit [1196:0] BITMAPS [43] = '{


        // <--- FILE: ASSETS\TEXT\REMATCH\REMATCH.PNG --->

        //tile 0, VRAM 48'b000000000000000000000000000001111101010100000000
        1197'b000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001000000001001001001001001001001001001001001001000000000001001001001001001001001001001001001001001001000000000001001001001001001001001001001001000000000000001001001001001001001001001001001001000000000000000000000000000001001001001001001001001001001001001000000000000001001001001001001001001001001001001000000001001001001001001000000000001001001001001001000001001001001001001001001001001001001001000001001001001001001000001001001001001001000000000001001001001001001000001001001001001001000000000001001001001001001000001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001000000001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001000000001001001001001001001001001001001001001001001000001001001001001001000000000001001001001001001000000000001001001001001001001001001001001000000000001001001001001001001001001001001001001000000000001001001001001001001001001001001000000000001001001001001001000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000001010010010010010010010010010010010010001000000001010010010010010010010010010010010001000000000001010010010010010010010010010010010010010001000000000001010010010010010010010010010001000000000000001010010010010010010010010010010001000000000000000000000000000001010010010010010010010010010010001000000000000001010010010010010010010010010010001000000001010010010010001000000000001010010010010001000001010010010010010010010010010010010001001001010010010010001000001010010010010001000000000001010010010010001000001010010010010001000000000001010010010010001001001010010010010010010010010010010010010010001000000000000000000001010010010010010010010010010010010001000000001010010010010010010010010010010001000000000000000000000001010010010010010010010010010010010010001000000001010010010010010010010010010010010010010001001001010010010010001000000000001010010010010001000000000001010010010010010010010010010001000000000001010010010010010010010010010010010001000000000001010010010010010010010010010001000000000001010010010010001000000001010010010010010001000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000001010010010010010010010010010010010010001001000001010010010010010010010010010010010001001001000001010010010010010010010010010010010010010001001001001001010010010010010010010010010001001001000001001010010010010010010010010010010001001001000000000000000001001001010010010010010010010010010010001001000001001001010010010010010010010010010010001001000001010010010010001001001001001010010010010001001001010010010010010010010010010010010001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001001000000000000000001010010010010010010010010010010010001001001001010010010010010010010010010010001001001000000000000000001010010010010010010010010010010010010001001000001010010010010010010010010010010010010010001001001010010010010001001001001001010010010010001001001001001010010010010010010010010010001001001000001010010010010010010010010010010010001001001001001010010010010010010010010010001001001000001010010010010001001001001010010010010010001001000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001001001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001000000000000000001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001000001010010010010010010001001001010010010010001001001010010010010010010010010010010010001001001010010010010001001001010010010010010010001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001001000000000000000001010010010010010010010010010010010001001001010010010010010010010010010010010010010001000000000000000001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001001001010010010010010010001010010010010010010001001001001010010010010010010010010010010010010001000001010010010010010010010010010010010001001001010010010010010010010010010010010010010001000001010010010010001001001001010010010010010001001000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000001010010010010010001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001001010010010010001001001001001010010010010001001001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010010001001001001010010010010001001001010010010010010010001001001010010010010001001001001001001010010010010010001001001001001001010010010010001001001010010010010010010001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001000000000000000001001001001010010010010001001001001001001001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010001001001001001001001001001001001001010010010010010010001010010010010010010001001001010010010010001001001001001010010010010001001001001001001010010010010001001001001001001001010010010010001001001001001010010010010001001001010010010010001001001001010010010010010001001000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000001010010010010010001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001001010010010010001001001001001010010010010001001001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010010001001001001010010010010001001001010010010010010010010010001010010010010001001001000000001010010010010010001001001001001001010010010010001001001010010010010010010010010001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001000000000000000000000000001010010010010001001001001001001001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010001001001001001001001001001001001001010010010010010010010010010010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010001001001001001001001010010010010001001001001001010010010010001001001010010010010001001001001010010010010010001001000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000001010010010010010001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001001010010010010001001001001001001001001001001001001010010010010001001001001001001001001001001001000000000000001010010010010010001001001001001001001001001001001010010010010010001001001001010010010010001001001010010010010010010010010001010010010010001001001000000001010010010010010001001001001001001010010010010001001001010010010010010010010010001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001000000000000000000000000001010010010010001001001001001001001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010001001001001001001001001001001001001010010010010010010010010010010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010001001001001001001001010010010010001001001001001001001001001001001001010010010010001001001001010010010010010001001000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000001010010010010010001001001001010010010010001001001010010010010010010010010010010010001001001001001010010010010010010010010010010010001001001000001001001010010010010010010010010010001001001001001001010010010010010010010010010010001001001001000000000000001010010010010010001001001001001001001001001001001010010010010010001001001001010010010010001001001010010010010001010010010010010010010010001001001000000001010010010010010001001000000000001010010010010001001001010010010010001010010010010010010010010001001001010010010010001001001001001010010010010001001001010010010010010010010010010010010001001001000000000000000000000000000001010010010010001001001000000000001010010010010001001001001010010010010010001001000000000000001010010010010010010010010010010010010001001001001010010010010010010010010010010010001001001000001010010010010001010010010001010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010001001001000000000001010010010010001001001001001001001001001001001001010010010010010010010010010010010010010001001000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000001010010010010010010010010010010010010010001001001010010010010010010010010010010010010010001001001010010010010010010010010010010010001001001000001001001010010010010010010010010010010010001001001001010010010010010010010010010010010010001001000000000000001010010010010010001001001001001001001001001001001010010010010010001001001001010010010010001001001010010010010001010010010010010010010010001001001000000001010010010010010001001000000000001010010010010001001001010010010010001010010010010010010010010001001001010010010010001001001001001010010010010001001001010010010010010010010010010010010001001001000000000000000000000000000001010010010010001001001000000000001010010010010001001001001010010010010010001001000000000000001010010010010010010010010010010010010010001001001010010010010010010010010010010010001001001000001010010010010001010010010001010010010010001001001010010010010010010010010010010010010010001001001000000001010010010010001001001000000000001010010010010001001001001001001001001001001000001010010010010010010010010010010010010010001001000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000001010010010010010010010010010010010010001001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001000001001001001001001001001001001010010010010001001001001001001001001001001001010010010010010001001000000000000001010010010010010001001001001001001001001001000001010010010010010001001001001010010010010001001001010010010010001001001010010010010010010001001001000000001010010010010010001001000000000001010010010010001001001010010010010001001001010010010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001000000000000000000000000000001010010010010001001001000000000001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010001001001001001001001001001001000001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001001001000000001010010010010001001001000000000001010010010010001001001001001001001001001001000001010010010010001001001001010010010010010001001000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000001010010010010010010010010010010010010001001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001000001010010010010001001001001001010010010010001001001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001000001010010010010010001001001001010010010010001001001010010010010001001001010010010010010010001001001000000001010010010010010001001000000000001010010010010001001001010010010010001001001010010010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001000000000000000000000000000001010010010010001001001000000000001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010001001001001001001001001001001000001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001001001000000001010010010010001001001000000000001010010010010001001001001001010010010010001000001010010010010001001001001010010010010010001001000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000001010010010010010001001001001001001001001001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001000001010010010010001001001001001010010010010001001001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010010001001001001010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010010001001000000000001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001000000000000000000000000000001010010010010001001001000000000001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010001001001001001001001001001001000001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010001001001000000000001010010010010001001001001001010010010010001001001010010010010001001001001010010010010010001001000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000001010010010010010001001001001001001001001001000001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001001001010010010010010010010010010010010010010001001000000000000001010010010010010010010010010010010010010001001001010010010010010010010010010010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010010001001000000000001010010010010001001001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001001001010010010010010010010010010010010010010001000000000000000000000000000001010010010010001001001000000000001010010010010010010010010010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010010010010010010010010010010001000001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010001001001000000000001010010010010010010010010010010010010010001001001010010010010001001001001010010010010010001001000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000001010010010010010001001001001001001001001001000001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001001001001001010010010010010010010010010001001001001001001010010010010010010010010010010001001001001000000000000001001001010010010010010010010010010010001001001001001001010010010010010010010010010010001001001001010010010010001001001001001010010010010001001001000000001010010010010010001001000000000001010010010010001001001010010010010001001001001001010010010010001001001001001010010010010010010010010010001001001001001010010010010010010010010010010010010010001001000000000000000000000000001010010010010001001001000000000001001010010010010010010010010010010001001001001000000000000001010010010010010001001001001010010010010001001001010010010010010010010010010010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001000000001010010010010001001001000000000001001001010010010010010010010010010001001001001001010010010010001001001001010010010010010001001000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000001001001001001001001001000000000001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000001001001001001001001001000000000000001001001001001001001001001001001001001001001000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000001001001001001001001001000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000001001001001001001000000000001001001001001001001001001001001001001001001001001001001001001001000000001001001001001001001001001001001001000000000000001001001001001001001001001001001001000000000000000000000000000001001001001001001001001001001001000000000000000001001001001001001001001001001001000000001001001001001001001000000000001001001001001001000000000000001001001001001001000000000000000001001001001001001000001001001001001001000000000001001001001001001000000001001001001001001001001001001001001000000001001001001001001001001001001001001001001001000000000000000000000000000000001001001001001001000000000000000000001001001001001001001001001001001001000000000000000000000001001001001001001000000000001001001001001001000001001001001001001001001001001001001001001001000001001001001001001000000000001001001001001001001001001001001001001000000001001001001001001001000000000000001001001001001001000000000000000000001001001001001001001001001001001001000000001001001001001001001000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000001001001001001001000000000001001001001001001000001001001001001001001001001001001001001001001000000001001001001001001001001001001001001000000000000001001001001001001001001001001001001000000000000000000000000000001001001001001001001001001001001000000000000000001001001001001001001001001001001000000000001001001001001001000000000001001001001001001000000000000001001001001001001000000000000000001001001001001001000001001001001001001000000000001001001001001001000000001001001001001001001001001001001001000000001001001001001001001001001001001001001001001000000000000000000000000000000001001001001001001000000000000000000001001001001001001001001001001001001000000000000000000000001001001001001001000000000001001001001001001000001001001001001001001001001001001001001001001000001001001001001001000000000001001001001001001000001001001001001001000000001001001001001001001000000000000001001001001001001000000000000000000001001001001001001001001001001001001000000001001001001001001001000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        1197'b001001001001001001001001001001001001001000000000001001001001001001001001001001001001001000000000001001001001001001001001001001001001001001001000000001001001001001001001001001001001001000000000000001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001000000000001001001001001001001001001001001001001001001000000001001001001001001001001001001001001000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000001001001001001001001001001001001001001001000000001001001001001001001001001001001001000000000000000000000001001001001001001001001001001001001001001000000001001001001001001001001001001001001001001001000001001001001001001001001001001001001001000001001001001001001000000000001001001001001001000001001001001001001001001001001001001001000000000001001001001001001000000000001001001001001001000000000000000000001001001001001001001001001001001001001000000001001001001001001001001001001001001000000000000000000000001001001001001001001000000001001001001001001000001001001001001001001001001001001001001001001000001001001001001001000000000001001001001001001000001001001001001001000000000001001001001001001000000,
        1197'b001010010010010010010010010010010010001000000000001010010010010010010010010010010010001000000000001010010010010010010010010010010010010010001000000001010010010010010010010010010010001000000000000001010010010010010010010010010010001000000000000000000000001010010010010010010010010010010010001000000000001010010010010010010010010010010010010010001000000001010010010010010010010010010010001000000000001010010010010010010010010010010010010010001001010010010010010010010010010010010010001000000000000000001010010010010010010010010010010010010001000000001010010010010010010010010010010001000000000000000000000001010010010010010010010010010010010010001000000001010010010010010010010010010010010010010001001001010010010010010010010010010010010001000001010010010010001000000000001010010010010001000001010010010010010010010010010010010001000000000001010010010010001000000000001010010010010001000000000000000000001010010010010010010010010010010010001000000001010010010010010010010010010010001000000000000000000000001010010010010010001000000001010010010010001000001010010010010010010010010010010010010010001000001010010010010001000000000001010010010010001000001010010010010001000000000001010010010010001000000,
        1197'b001010010010010010010010010010010010001001001000001010010010010010010010010010010010001001001000001010010010010010010010010010010010010010001001001001010010010010010010010010010010001001000001001001010010010010010010010010010010001001000000000000000000001010010010010010010010010010010010001001001000001010010010010010010010010010010010010010001001001001010010010010010010010010010010001001001000001010010010010010010010010010010010010010001001010010010010010010010010010010010010001001000000000000001010010010010010010010010010010010010001001001001010010010010010010010010010010001001001000000000000000001010010010010010010010010010010010010001001000001010010010010010010010010010010010010010001001001010010010010010010010010010010010001001001010010010010001001001001001010010010010001001001010010010010010010010010010010010001001001000001010010010010001001001001001010010010010001001001000000000000001010010010010010010010010010010010001001001001010010010010010010010010010010001001001000000000000000001010010010010010001001001001010010010010001001001010010010010010010010010010010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001,
        1197'b001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001000000000000000000001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001001001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001001010010010010010010010010010010010010001001000000000000001010010010010010010010010010010010010001001001010010010010010010010010010010010010010001000000000000000001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001001001010010010010010010010010010010010001001001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001000001010010010010010010001001001010010010010001001001000000000000001010010010010010010010010010010010001001001010010010010010010010010010010010010010001000000000000000001010010010010010010001010010010010010010001001001010010010010010010010010010010010010010001001001010010010010010010001001001010010010010001001001010010010010001001001001001010010010010001001001,
        1197'b001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001010010010010010001001001001010010010010001001001010010010010010001001001001010010010010001001001000000000000001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001001010010010010001001001001010010010010010001001001010010010010001001001001001001001001001001001001001001001010010010010001001001001001001000000000000001001001001001010010010010001001001001001001001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010001001001001001001001001001001001001001001001001010010010010001001001001001001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010010010001001001010010010010001001001000000000000001001001001010010010010001001001001001001001010010010010001001001001010010010010010001001000000000000001010010010010010010001010010010010010010001001001010010010010010001001001001001001001001001001001010010010010010010001001001010010010010001001001010010010010001001001001001010010010010001001001,
        1197'b001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001010010010010010001001001001010010010010001001001010010010010010001001001001010010010010001001001000000000000001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001001010010010010001001001001010010010010010001001001010010010010001001001001001001001001001001001000000000001010010010010001001001001001001000000000000000000000000001010010010010001001001001001001001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010001001001001001001001001001001001001000000000001010010010010001001001001001001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010010010010010001010010010010001001001000000000000000000000001010010010010001001001001001001001010010010010001001001001010010010010010001001000000000000001010010010010010010010010010010010010010001001001010010010010010001001001001001001001001001001001010010010010010010010010001010010010010001001001010010010010001001001001001010010010010001001001,
        1197'b001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001010010010010010001001001001001001001001001001001010010010010010001001001001001001001001001001001000000000000001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001001010010010010001001001001001001001001001001001001010010010010001001001001001001001001001001001000000000001010010010010001001001001001001000000000000000000000000001010010010010001001001001001001001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010001001001001001001001001001001001001000000000001010010010010001001001001001001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010010010010010001010010010010001001001000000000000000000000001010010010010001001001001001001001010010010010001001001001010010010010010001001000000000000001010010010010010010010010010010010010010001001001010010010010010001001001001001001001001001001001010010010010010010010010001010010010010001001001010010010010001001001001001010010010010001001001,
        1197'b001010010010010001001001001001010010010010001001001010010010010010010010010010010010001001001001001010010010010010010010010010010010001001001001001001010010010010010010010010010010001001001001001001010010010010010010010010010010001001001001000000000000001010010010010010010010010010010010001001001001001010010010010010010010010010010010001001001000001001010010010010010010010010010010001001001001001010010010010010010010010010010010001001001000000000000001010010010010001001001000000000000000000000000000000000001010010010010001001001000000000001010010010010001001001001010010010010010001001000000000000001010010010010010010010010010010010010001001001001010010010010010010010010010010010001001001000000000000000001010010010010001001001000000001010010010010001001001001001010010010010001001001010010010010010010010010010010010001001001001001010010010010001010010010010010010010010001001001000000000000000000000001010010010010001001001000000000001010010010010001001001001010010010010010001001000000000000001010010010010010001010010001010010010010001001001010010010010010010010010010010010010001001000001010010010010001010010010010010010010010001001001010010010010001001001001001010010010010001001001,
        1197'b001010010010010010010010010010010010010010001001001010010010010010010010010010010010010010001001001010010010010010010010010010010010001001001001001001010010010010010010010010010010010001001001001001010010010010010010010010010010010001001001000000000000001010010010010010010010010010010010010010001001001010010010010010010010010010010010001001001000001001010010010010010010010010010010010010001001001010010010010010010010010010010010001001001000000000000001010010010010001001001000000000000000000000000000000000001010010010010001001001000000000001010010010010001001001001010010010010010001001000000000000001010010010010010010010010010010010010010001001001010010010010010010010010010010010001001001000000000000000001010010010010001001001000000001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001001001010010010010001010010010010010010010010001001001000000000000000000000001010010010010001001001000000000001010010010010001001001001010010010010010001001000000000000001010010010010010001010010001010010010010001001001010010010010010010010010010010010010001001000001010010010010001010010010010010010010010001001001010010010010001001001001001010010010010001001001,
        1197'b001010010010010010010010010010010010001001001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001001001001001001001001001001010010010010001001001001001001001001001001001001010010010010001001001000000000000001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001000001001001001001001001001001010010010010010001001001010010010010001001001001001001001001001001000000000000001010010010010001001001000000000000000000000000000000000001010010010010001001001000000000001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010001001001001001001001001001001000000000000000001010010010010001001001000000001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001010010010010010010001001001000000000000000000000001010010010010001001001000000000001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010010001001001001001001001001001000001010010010010001001001010010010010010010001001001010010010010001001001001001010010010010001001001,
        1197'b001010010010010010010010010010010010001001001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001010010010010010001001001001010010010010001001001010010010010010001001001001010010010010001001001000000000000001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001000001010010010010001001001001010010010010010001001001010010010010001001001001001001001001001001000000000000001010010010010001001001000000000000000000000000000000000001010010010010001001001000000000001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010001001001001001001001001001001000000000000000001010010010010001001001000000001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001010010010010010010001001001000000000000000000000001010010010010001001001000000000001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010010001001001001001001001001001000001010010010010001001001010010010010010010001001001010010010010001001001001001010010010010001001001,
        1197'b001010010010010001001001001001001001001001001001001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001001010010010010010001001001001010010010010001001001010010010010010001001001001010010010010001001001000000000000001010010010010001001001001001010010010010001001001010010010010001001001001001001001001001001000001010010010010001001001001010010010010010001001001010010010010001001001001001001001001001001000000000000001010010010010001001001000000000000000000000000000000000001010010010010001001001000000000001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010001001001001001001001001001001000000000000000001010010010010001001001000000001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001000000000000000000000001010010010010001001001000000000001010010010010001001001001010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010010001001001001001001001001001000001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001,
        1197'b001010010010010001001001001001001001001001001000001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001001010010010010010010010010010010010010010001001001010010010010010010010010010010010010010001001001000000000000001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001000001010010010010010010010010010010010010010001001001010010010010010010010010010010010010010001000000000000001010010010010001001001000000000000000000000000000000000001010010010010001001001000000000001010010010010010010010010010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010010010010010010010010010010001000000000000000001010010010010001001001000000001010010010010010010010010010010010010010001001001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001000000000000000000000001010010010010001001001000000000001010010010010010010010010010010010010010001001000000000000001010010010010010001001001001010010010010001001001010010010010010010010010010010010010010001001001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001001001,
        1197'b001010010010010001001001001001001001001001001000001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001001001001010010010010010010010010010010001001001001001001010010010010010010010010010010001001001001000000000000001010010010010001001001001001010010010010001001001010010010010010010010010010010010010010001001001001010010010010010010010010010010001001001001001010010010010010010010010010010010010010001001000000000001010010010010001001001000000000000000000000000000000000001010010010010001001001000000000001001010010010010010010010010010010001001001001000000000000001010010010010010001001001001010010010010001001001010010010010010010010010010010010010010001001001000000000001010010010010001001001000000001001001010010010010010010010010010001001001001001010010010010001001001001001010010010010001001001010010010010001001001001001010010010010001001001000000000000000000000001010010010010001001001000000000001001010010010010010010010010010010001001001001000000000000001010010010010010001001001001010010010010001001001010010010010010010010010010010010010010001001001010010010010001001001001001010010010010001001001001001010010010010010010010010010001001001001001,
        1197'b001001001001001001001001000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000001001001001001001001001000000000000000000000000000000000001001001001001001001001000000000000001001001001001001001001001001001001001001001000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000001001001001001001001001000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000001001001001001001001001000000000000001001001001001001001001001001001001001001001000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000001001001001001001001001001001001001001001001,
        1197'b000000001001001001001001000000000000000000000000000000001001001001001001000000001001001001001001001001001001001001001001001001001001001001001001000000000001001001001001001001001001001001000000000000000001001001001001001001001001001001000000000000000000000000001001001001001001000000000001001001001001001001001001001001001001001001001001001001001001001000000001001001001001001001001001001001001000000001001001001001001001001001001001001001001001000000000000000001001001001001001000000000000000000000000000000000000000001001001001001001000000000000000000001001001001001001001001001001001001000000000000000000000001001001001001001000000000001001001001001001000001001001001001001001001001001001001001001001000000000000001001001001001001001000000000000000000001001001001001001001001001001001001000000001001001001001001000000001001001001001001001001001001001001001001000000001001001001001001001000000000000000000000000000001001001001001001000000000000000000001001001001001001001001001001001001000000000000000000000001001001001001001000000000001001001001001001000001001001001001001001001001001001001001001001000001001001001001001000000000001001001001001001000000001001001001001001001001001001001001000000,
        1197'b000000001001001001001001000000000000000000000000000000001001001001001001000000001001001001001001001001001001001001001001001001001001001001001001000000000001001001001001001001001001001001000000000000000001001001001001001001001001001001000000000000000000000000001001001001001001000000000001001001001001001000001001001001001001001001001001001001001001001000000001001001001001001001001001001001001000000001001001001001001001001001001001001001001001000000000000000001001001001001001000000000000000000000000000000000000000001001001001001001000000000000000000001001001001001001001001001001001001000000000000000000000001001001001001001000000000001001001001001001000001001001001001001001001001001001001001001001000000000000001001001001001001001000000000000000000001001001001001001001001001001001000000000001001001001001001000000001001001001001001001000001001001001001001000000001001001001001001001000000000000000000000000000001001001001001001000000000000000000001001001001001001001001001001001001000000000000000000000001001001001001001000000000001001001001001001000001001001001001001001001001001001001001001001000001001001001001001000000000001001001001001001000000001001001001001001001001001001001001000000
    
    };

    always_comb
    begin
        bitmapIdx = PixelY;
        bitmap    = BITMAPS[bitmapIdx];
        color     = bitmap[3*(398-PixelX) +: 3];
        Data      = data[6*color+0 +: 6];
    end

endmodule
