module money_rom (
    input  logic [1:0]  Tile,
    input  logic [4:0] PixelX,
    input  logic [4:0] PixelY,
    output logic [5:0]  Data
);

    logic [49:0] data;
    logic [6:0] bitmapIdx;
    logic [77:0] bitmap;
    logic [2:0]  color;

    localparam bit [49:0] DATA [3] = '{


        // <--- FILE: MONEY\PALLETS.PNG --->

        //tile 0
        50'b00000000000000000001100110110100010010110000000000,
        //tile 1
        50'b00111001100110111010110100010000111110110000000001,
        //tile 2
        50'b11000001100110111110111010110100010010110000000010
    
    };

    localparam bit [77:0] BITMAPS [84] = '{


        // <--- FILE: MONEY\PALLETS.PNG --->

        //tile 0, VRAM 50'b00000000000000000001100110110100010010110000000000
        78'b000000000001001001001000000001001001001000000001001001001000000001001001001000,
        78'b000000010001001001001000010001001001001000010001001001001000010001001001001000,
        78'b000011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b000011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b010011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b010011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b010100100001001001001100100001001001001100100001001001001100100001001001001100,
        78'b010010010001001001001010010001001001001010010001001001001010010001001001001000,
        78'b000011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b000011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b010011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b010011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b010100100001001001001100100001001001001100100001001001001100100001001001001100,
        78'b010010010001001001001010010001001001001010010001001001001010010001001001001000,
        78'b000011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b000011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b010011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b010011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b010100100001001001001100100001001001001100100001001001001100100001001001001100,
        78'b010010010001001001001010010001001001001010010001001001001010010001001001001000,
        78'b000011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b000011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b010011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b010011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b010100100001001001001100100001001001001100100001001001001100100001001001001100,
        78'b010010010001001001001010010001001001001010010001001001001010010001001001001000,
        78'b000000010011011011011000010011011011011000010011011011011000010011011011011000,
        78'b000000010010010010000000010010010010000000010010010010000000010010010010000000,
        //tile 1, VRAM 50'b00111001100110111010110100010000111110110000000001
        78'b000000000001001001001010010010010010010000010010010010010010000001001001001000,
        78'b000000011001010010010010011010010011010010010011010010011010010010010010001000,
        78'b000100100001010011010010010010010010010010010010010010010010010010011010001100,
        78'b000100100001010010010010010010010010010010010010010010010010010010010010001100,
        78'b011100100001010010010101101101101101101010101101101101101101010010010010001100,
        78'b011100100001101101101101101101101010010010010010010101101101101101101101001100,
        78'b011110110001101101101010010010010010011010010011010010010010101101101101001110,
        78'b011011011001010010010010010010010010010010010010010010010010010010010010001000,
        78'b000100100001010010010010011010010010010010010010010010011010010010010010001100,
        78'b000100100001010011010010010010010101101101101101101010010010010010011010001100,
        78'b011100100001010010010111111111111101101101101101101111111111010010010010001100,
        78'b011100100001111111111010010010010010010010010010010010010010111111111111001100,
        78'b011110110001001001001010011010010010010010010010010010011010110001001001001110,
        78'b011011011001010010010010010010010010011010010011010010010010010010010010001000,
        78'b000100100001010011010010010010010010010010010010010010010010010010011010001100,
        78'b000100100001010010010101101101101111111111111111111101101101010010010010001100,
        78'b011100100001010010010101101101101101101010101101101101101101010010010010001100,
        78'b011100100001101101101010010010010010010101010010010010010010101101101101001100,
        78'b011110110001101101101010010010010010010101010010010010010010101101101101001110,
        78'b011011011001010010010010011010010011010010010011010010011010010010010010001000,
        78'b000100100001010010010010010010010010010010010010010010010010010010010010001100,
        78'b000100100001010011010111111111111111111010111111111111111111010010011010001100,
        78'b011100100001010010010010010010001010010010010010010001010010010010010010001100,
        78'b011100100001111111111111111111001111111111111111111001111111111111111111001100,
        78'b011110110001001001001110110001001001001110110001001001001110110001001001001110,
        78'b011011011001001001001011011001001001001011011001001001001011011001001001001000,
        78'b000000011100100100100000011100100100100000011100100100100000011100100100100000,
        78'b000000011011011011000000011011011011000000011011011011000000011011011011000000,
        //tile 2, VRAM 50'b11000001100110111110111010110100010010110000000010
        78'b000000000001001001001000000001001001001000000001001001001000000001001001001000,
        78'b000000010001001001001000010001001001001000010001001001001000010001001001001000,
        78'b000011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b000011011001001100100011011100100001001100100001001100100011011100100001001011,
        78'b010011011001101100100101101100100101101100100101101100100101101100100101001011,
        78'b010011011001101100100101101100100101101100100101101100100101101100100101001011,
        78'b010110110001101100100101101100100101101100100101101100100101101100100101100110,
        78'b010010010001101100100101101100100101101100100101101100100101101100100101100000,
        78'b000011011001101100100101101100100101101100100101101100100101101100100101100011,
        78'b000011011001101100100101101100100101101100100101101100100101101100100101100011,
        78'b010011011001101111111101101111111101101111111101101111111101101111111101100011,
        78'b010011011001100100111111100100111111100100111111100100111111100100111111100011,
        78'b010110110101100100101101100100101101100100101101100100101101100100101111100110,
        78'b010010010101100100101101100100101101100100101101100100101101100100101111111000,
        78'b000011011101100100101101100100101101100100101101100100101101100100101100001011,
        78'b000011011101100100101101100100101101100100101101100100101101100100101100001011,
        78'b010011011101100100101101100100101101100100101101100100101101100100101100001011,
        78'b010011011101100100101101100100101101100100101101100100101101100100101100001011,
        78'b010110110101111111101101111111101101111111101101111111101101111111101100001110,
        78'b010010010111111111111111111111111111111111111111111111111111111111111100001000,
        78'b000011011101101111111101101111111101101111111101101111111101101111111100001011,
        78'b000011011101111111111111111111111111111111111111111111111111111111111111001011,
        78'b010011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b010011011001001001001011011001001001001011011001001001001011011001001001001011,
        78'b010110110001001001001110110001001001001110110001001001001110110001001001001110,
        78'b010010010001001001001010010001001001001010010001001001001010010001001001001000,
        78'b000000010011011011011000010011011011011000010011011011011000010011011011011000,
        78'b000000010010010010000000010010010010000000010010010010000000010010010010000000
    
    };

    always_comb
    begin
        data      = DATA[Tile];
        bitmapIdx = 28 * data[1:0] + PixelY;
        bitmap    = BITMAPS[bitmapIdx];
        color     = bitmap[3*(25-PixelX) +: 3];
        Data      = data[6*color+2 +: 6];
    end

endmodule
