module map_rom (
    input  logic [10:0]  Tile,
    input  logic [3:0] PixelX,
    input  logic [3:0] PixelY,
    output logic [5:0]  Data
);

    logic [55:0] data;
    logic [11:0] bitmapIdx;
    logic [47:0] bitmap;
    logic [2:0]  color;

    localparam bit [55:0] DATA [1200] = '{


        // <--- FILE: MAP\CITY.PNG --->

        //tile 0
        56'b00000000000000000000000000010000001100001000000100000000,
        //tile 1
        56'b00000000000000000000000000010000001100001000000100000000,
        //tile 2
        56'b00000000000000000000000000010000001100001000000100000000,
        //tile 3
        56'b00000000000000000000000000010000001100001000000100000000,
        //tile 4
        56'b00000000000000000000000000001100010000001000000100000001,
        //tile 5
        56'b00000000000000000000100100100000011100011000010100000010,
        //tile 6
        56'b00000000000000000000000000100100100000010100011000000011,
        //tile 7
        56'b00000000000000000000000000100100100000010100011000000011,
        //tile 8
        56'b00000000000000000000100100100000011100010100011000000100,
        //tile 9
        56'b00000000000000000000001000101000001100000100010000000101,
        //tile 10
        56'b00000000000000000000001000010000001100000100101000000110,
        //tile 11
        56'b00000000000000000000001000010000001100000100101000000110,
        //tile 12
        56'b00000000000000000000001000010000001100000100101000000111,
        //tile 13
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 14
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 15
        56'b00000000001000001100110100110000101100010000000100001001,
        //tile 16
        56'b00000000000000000000000000001000001100000100010000001010,
        //tile 17
        56'b00000001001001000101000000111100101000010000111000001011,
        //tile 18
        56'b00000000000000000000000001001100111100111000010000001100,
        //tile 19
        56'b00000000000000000000000000000001001100111000111100001101,
        //tile 20
        56'b00000000000000000000000000010000111001001100111100001110,
        //tile 21
        56'b00000000000000000000000000001000001100000100010000001010,
        //tile 22
        56'b00000000001000001100000100101100110000110100010000001111,
        //tile 23
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 24
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 25
        56'b00000000000000000000100100100000011100011000010100000010,
        //tile 26
        56'b00000000000000000000000000100100100000010100011000000011,
        //tile 27
        56'b00000000000000000000000000100100100000010100011000000011,
        //tile 28
        56'b00000000000000000000000000100100100000010100011000000011,
        //tile 29
        56'b00000000000000000000000000100100100000010100011000000011,
        //tile 30
        56'b00000000000000000000100100100000011100010100011000000100,
        //tile 31
        56'b00000000000000000000000001011101011001010101010000010000,
        //tile 32
        56'b00000000000000000000000001011101011001010101010000010001,
        //tile 33
        56'b00000000000000000000000001011101011001010101010000010001,
        //tile 34
        56'b00000000000000000000000001011101011001010101010000010001,
        //tile 35
        56'b00000000000000000000000001011101011001010101010000010001,
        //tile 36
        56'b00000000000000000000000001011101011001010101010000010010,
        //tile 37
        56'b00000000000000000000000001101101101001100101100000010011,
        //tile 38
        56'b00000000000000000000000001100001101101101001100100010100,
        //tile 39
        56'b00000000000000000000000001101101101001100001100100010101,
        //tile 40
        56'b00000000000000000000000000101000001100000100001000010110,
        //tile 41
        56'b00000000000000000000000000101000001100000100001000010110,
        //tile 42
        56'b00000000000000000000000000101000001100000100001000010110,
        //tile 43
        56'b00000000000000000000000000101000001100000100001000010110,
        //tile 44
        56'b00000000000000000000000000101000001100000100001000010111,
        //tile 45
        56'b00000000000000000000000000000001101101100001100100011000,
        //tile 46
        56'b00000000000000000000000000000001100101101101100000011001,
        //tile 47
        56'b00000000000000000000000000000001100101101101100000011001,
        //tile 48
        56'b00000000000000000000000000000001101101100101100000011010,
        //tile 49
        56'b00000000000000000000000001010101010001011101110000011011,
        //tile 50
        56'b00000000000000000000000001010101010001110001011100011100,
        //tile 51
        56'b00000000000000000000000001010101010001110001011100011100,
        //tile 52
        56'b00000000000000000000000001010101010001110001011100011101,
        //tile 53
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 54
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 55
        56'b00000000110000101100110100001100010000001000000100011110,
        //tile 56
        56'b00000000000000000000000000001000001100000100010000001010,
        //tile 57
        56'b00000001001001000101000000111100101000010000111000001011,
        //tile 58
        56'b00000001000001001001000100111101001100010000111000011111,
        //tile 59
        56'b00000000011100010101110000111100010000111001001100100000,
        //tile 60
        56'b00000000000001000000111100101000111000010001001100100001,
        //tile 61
        56'b00000000000000000000000000001000001100000100010000001010,
        //tile 62
        56'b00000000101100110000001100110100000100010000001000100010,
        //tile 63
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 64
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 65
        56'b00000000000000000000000000010100011100100101110100100011,
        //tile 66
        56'b00000000000000000000000000010100011101110100100100100100,
        //tile 67
        56'b00000000000000000000000000010100011101110100100100100100,
        //tile 68
        56'b00000000000000000000000000010100011101110100100100100100,
        //tile 69
        56'b00000000000000000000000000010100011101110100100100100100,
        //tile 70
        56'b00000000000000000000000000010100011101110100100100100101,
        //tile 71
        56'b00000000000000000000101001111000001100000100001000100110,
        //tile 72
        56'b00000000000000000000101001111000001100000100001000100111,
        //tile 73
        56'b00000000000000000000000000101000001100000100001000101000,
        //tile 74
        56'b00000000000000000000000000101000001100000100001000101001,
        //tile 75
        56'b00000000000000000000101001111000001100000100001000100111,
        //tile 76
        56'b00000000000000000000101001111000001100000100001000101010,
        //tile 77
        56'b00000000000000000000000000000001101101100001100100011000,
        //tile 78
        56'b00000000001100010000111000000100111100101000001000101011,
        //tile 79
        56'b00000000000000000000000000000001101101100101100000011010,
        //tile 80
        56'b00000000000000000000101001111000001100000100001000101100,
        //tile 81
        56'b00000000000000000000000000010000000100001001111000101101,
        //tile 82
        56'b00000000000000000000000000010000000100001001111000101110,
        //tile 83
        56'b00000000000000000000101001111000001100000100001000101111,
        //tile 84
        56'b00000000000000000000101001111000001100000100001000110000,
        //tile 85
        56'b00000000000000010000111000000100111100101000001000110001,
        //tile 86
        56'b00000000000000010000000100111000101000111100001000110010,
        //tile 87
        56'b00000000000000000001100001010001011001011101010100110011,
        //tile 88
        56'b00101100110000101000100001100001100100010000001000110100,
        //tile 89
        56'b00000000000000000000000001010101010001011101110000110101,
        //tile 90
        56'b00000000000000000000000000001000001100000100101000110110,
        //tile 91
        56'b00000000000000000000000000001000001100000100101000110110,
        //tile 92
        56'b00000000000000000000000001010101010001011101110000110101,
        //tile 93
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 94
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 95
        56'b00000000001000001100110100110000101100010000000100001001,
        //tile 96
        56'b00000000000000000000000000001000001100000100010000110111,
        //tile 97
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 98
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 99
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 100
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 101
        56'b00000000000000000000000000001000010000000100001100111001,
        //tile 102
        56'b00000000001000001100000100101100110000110100010000001111,
        //tile 103
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 104
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 105
        56'b01011001111100100101101000011101110100010000001000111010,
        //tile 106
        56'b01100001101101100100111000010000111100101000001000111011,
        //tile 107
        56'b01100001101101100100010000111000101000111100001000111100,
        //tile 108
        56'b00000001111000010000111000000100111100101000001000111101,
        //tile 109
        56'b00000001111000010000000100111000101000111100001000111110,
        //tile 110
        56'b00000000111001011101000001110100011100010000001000111111,
        //tile 111
        56'b00000000000000000000101001111000001100000100001000100110,
        //tile 112
        56'b00000000000000000000101001111000001100000100001000101010,
        //tile 113
        56'b00000000000000000000000000010000000100001001111000101101,
        //tile 114
        56'b00000000000000000000000000010000000100001001111000101110,
        //tile 115
        56'b00000000000000000000101001111000001100000100001000100110,
        //tile 116
        56'b00000000000000000000101001111000001100000100001000101010,
        //tile 117
        56'b01100001101101100100111000010000111100101000001001000000,
        //tile 118
        56'b00000100101001000100110101100101100000010000001001000001,
        //tile 119
        56'b00000000001100010000111000000100111100101000001000101011,
        //tile 120
        56'b00000000000000000000000000000000001100001000000101000010,
        //tile 121
        56'b00000000000000000000000000000100010000001001111001000011,
        //tile 122
        56'b00000000000000000000000000000100001000010001111001000100,
        //tile 123
        56'b00000000000000000000000000000000001100000100001001000101,
        //tile 124
        56'b00000000000000000000000000000000001100001000000101000010,
        //tile 125
        56'b00000000000000000000000000000001101101100001100100011000,
        //tile 126
        56'b00000000000000000000000000000001101101100101100000011010,
        //tile 127
        56'b00000001101001010001000001100001011001011101010101000110,
        //tile 128
        56'b00000000000000000000000000000001101101100001100101000111,
        //tile 129
        56'b00000000000000000000000001010101010001011101110000110101,
        //tile 130
        56'b00000000000000000000000000001000001100000100101000110110,
        //tile 131
        56'b00000000000000000000000000001000001100000100101000110110,
        //tile 132
        56'b00000000000000000000000001010101010001011101110000110101,
        //tile 133
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 134
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 135
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 136
        56'b00000000110000001100101100110100000100010000001001001000,
        //tile 137
        56'b00000000001100110000101100000100110100001000010001001001,
        //tile 138
        56'b00000000111001001100111100001100010000001000000101001010,
        //tile 139
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 140
        56'b00000000110000001100101100110100000100010000001001001000,
        //tile 141
        56'b00000000001100110000101100000100110100001000010001001001,
        //tile 142
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 143
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 144
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 145
        56'b00000000000000000000000000010100011100100101110101001011,
        //tile 146
        56'b00000000000000000000000000000001100001101101100101001100,
        //tile 147
        56'b00000000000000000000000000000001100001101101100101001101,
        //tile 148
        56'b00000000000000000000000000010100011100100101110100100011,
        //tile 149
        56'b00000000000000000000000000010100011101110100100100100100,
        //tile 150
        56'b00000000000000000000000000010100011101110100100100100101,
        //tile 151
        56'b00000000000000000000000000000000001100000100001001000101,
        //tile 152
        56'b00000000000000000000000000000000001100001000000101000010,
        //tile 153
        56'b00000000000000000000000000000100010000001001111001000011,
        //tile 154
        56'b00000000000000000000000000000100001000010001111001000100,
        //tile 155
        56'b00000000000000000000000000000000001100000100001001000101,
        //tile 156
        56'b00000000000000000000000000000000001100001000000101000010,
        //tile 157
        56'b00000000000000000000000000000001100001101101100101001100,
        //tile 158
        56'b00000000000000000000000000000001100101101101100000011001,
        //tile 159
        56'b00000000000000000000000000000001101101100101100000011010,
        //tile 160
        56'b00111000001100111101001110000000010000001000000101001110,
        //tile 161
        56'b00000000000000000000000000001000001100000100010001001111,
        //tile 162
        56'b00000000000000000000000000001000010000000100001101010000,
        //tile 163
        56'b00000000110000001100101100110100000100010000001001001000,
        //tile 164
        56'b00000000001100110000101100000100110100001000010001001001,
        //tile 165
        56'b00111000001100111101001110000000010000001000000101001110,
        //tile 166
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 167
        56'b00000000000000000000000000001000001100000100010001010001,
        //tile 168
        56'b00000000111001001100111100001100010000001000000101001010,
        //tile 169
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 170
        56'b00000000000000000000000000001000001100000100010001010010,
        //tile 171
        56'b00000000000000000000000000001000010000000100001101010011,
        //tile 172
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 173
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 174
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 175
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 176
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 177
        56'b00000010010010001110001010000100001100001000000101010100,
        //tile 178
        56'b00000000000010001010010110010010001110000100000101010101,
        //tile 179
        56'b00000000000000000000000000000010010010001110000101010110,
        //tile 180
        56'b00000000000000000000000010010010001100000110000101010111,
        //tile 181
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 182
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 183
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 184
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 185
        56'b00111000001100111101001110000000010000001000000101001110,
        //tile 186
        56'b00000000000000000000000000001000001100000100010001001111,
        //tile 187
        56'b00000000000000000000000000001000010000000100001101010000,
        //tile 188
        56'b00111000001100111101001110000000010000001000000101001110,
        //tile 189
        56'b00000000110000001100101100110100000100010000001001001000,
        //tile 190
        56'b00000000001100110000101100000100110100001000010001001001,
        //tile 191
        56'b00111000001100111101001110000000010000001000000101001110,
        //tile 192
        56'b00111000111100001101000000101000010000001000000101011000,
        //tile 193
        56'b00000000000000000000000000001000001100000100010001001111,
        //tile 194
        56'b00000000000000000000000000001000010000000100001101010000,
        //tile 195
        56'b00111000111100001101000000101000010000001000000101011000,
        //tile 196
        56'b00111000001100111101001110000000010000001000000101001110,
        //tile 197
        56'b00000000000000000000000000001000001100000100010001010001,
        //tile 198
        56'b00000000110000001100101100110100000100010000001001001000,
        //tile 199
        56'b00000000001100110000101100000100110100001000010001001001,
        //tile 200
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 201
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 202
        56'b00000000000000000000000000010000001100001000000101011001,
        //tile 203
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 204
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 205
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 206
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 207
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 208
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 209
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 210
        56'b00000000000000000000000000001000001100000100010001010010,
        //tile 211
        56'b00000000000000000000000000001000010000000100001101010011,
        //tile 212
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 213
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 214
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 215
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 216
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 217
        56'b00001000010000001100000110001010010010001110000101011010,
        //tile 218
        56'b00000000010010011010010010000110001110001010010101011011,
        //tile 219
        56'b00000000000000010000001010000110010010001010001101011100,
        //tile 220
        56'b00000000000000001000010000001110010010000110001101011101,
        //tile 221
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 222
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 223
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 224
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 225
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 226
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 227
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 228
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 229
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 230
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 231
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 232
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 233
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 234
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 235
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 236
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 237
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 238
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 239
        56'b00000000000000000000000000010000001100001000000101011001,
        //tile 240
        56'b00000001111101000001101000001100010000001000000101011110,
        //tile 241
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 242
        56'b00000000000000000000000000001100010000001000000101011111,
        //tile 243
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 244
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 245
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 246
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 247
        56'b00000001111101000001101000001100010000001000000101011110,
        //tile 248
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 249
        56'b00000000000000000000000000010000001100001000000101100000,
        //tile 250
        56'b00000000000000000000000000001000001100000100010001010010,
        //tile 251
        56'b00000000000000000000000000001000010000000100001101010011,
        //tile 252
        56'b00000000000000000000000000010000001100001000000101100000,
        //tile 253
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 254
        56'b00000001111101000001101000001100010000001000000101011110,
        //tile 255
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 256
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 257
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 258
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 259
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 260
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 261
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 262
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 263
        56'b00000001111101000001101000001100010000001000000101100001,
        //tile 264
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 265
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 266
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 267
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 268
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 269
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 270
        56'b00000001111101000001101000001100010000001000000101100001,
        //tile 271
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 272
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 273
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 274
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 275
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 276
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 277
        56'b00000001111101000001101000001100010000001000000101100001,
        //tile 278
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 279
        56'b00000000000000000000000000001100010000001000000101011111,
        //tile 280
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 281
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 282
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 283
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 284
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 285
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 286
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 287
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 288
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 289
        56'b00000000000000000000000000010000001100001000000101100011,
        //tile 290
        56'b00000000000000000000000000001000001100000100010001010010,
        //tile 291
        56'b00000000000000000000000000001000010000000100001101010011,
        //tile 292
        56'b00000000000000000000000000010000001100001000000101100011,
        //tile 293
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 294
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 295
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 296
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 297
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 298
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 299
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 300
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 301
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 302
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 303
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 304
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 305
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 306
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 307
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 308
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 309
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 310
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 311
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 312
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 313
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 314
        56'b00010001011100101001011000001101010100001000000101100100,
        //tile 315
        56'b00000000000000000001100000001101100100001000000101100101,
        //tile 316
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 317
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 318
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 319
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 320
        56'b00000000000000000000000000001000000100001100010001100110,
        //tile 321
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 322
        56'b00000000000000000000000000001000000100001100010001100110,
        //tile 323
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 324
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 325
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 326
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 327
        56'b00000000000000000000000000001000000100001100010001100111,
        //tile 328
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 329
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 330
        56'b00000000000000000000000000001000001100000100010001001111,
        //tile 331
        56'b00000000000000000000000000001000010000000100001101010000,
        //tile 332
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 333
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 334
        56'b00000000000000000000000000001000000100001100010001100111,
        //tile 335
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 336
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 337
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 338
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 339
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 340
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 341
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 342
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 343
        56'b00000000000000000000000000001000000100001100010001101000,
        //tile 344
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 345
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 346
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 347
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 348
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 349
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 350
        56'b00000000000000000000000000001000000100001100010001101000,
        //tile 351
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 352
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 353
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 354
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 355
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 356
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 357
        56'b00000000000000000000000000001000000100001100010001101001,
        //tile 358
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 359
        56'b00000000000000000000000000001000000100001100010001101010,
        //tile 360
        56'b00000000000000000000000000001000001100000100010001101011,
        //tile 361
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 362
        56'b00000000000000000000000000001000000100001100010001101100,
        //tile 363
        56'b00000000000000000000000000000000101000001000010001101101,
        //tile 364
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 365
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 366
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 367
        56'b00000000000000000000000000000000101000010000001001110000,
        //tile 368
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 369
        56'b00000000000000000000000000000000000000101000001001110001,
        //tile 370
        56'b00000000000000000000000000000000000000101000001001110001,
        //tile 371
        56'b00000000000000000000000000000000000000101000001001110001,
        //tile 372
        56'b00000000000000000000000000000000000000101000001001110001,
        //tile 373
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 374
        56'b00000000000000000000000000000000101000010000001001110010,
        //tile 375
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 376
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 377
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 378
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 379
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 380
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 381
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 382
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 383
        56'b00000000000000000000000000000000101000010000001001110011,
        //tile 384
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 385
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 386
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 387
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 388
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 389
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 390
        56'b00000000000000000000000000000000101000010000001001110100,
        //tile 391
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 392
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 393
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 394
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 395
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 396
        56'b00000000000000000000000000000000000000101000001001110101,
        //tile 397
        56'b00000000000000000000000000001000001100000100010001110110,
        //tile 398
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 399
        56'b00000000000000000000000000001000000100001100010001101100,
        //tile 400
        56'b00000000000000000000000000000000000000101000001001110111,
        //tile 401
        56'b00000000000000000000000000000000000000001000101001111000,
        //tile 402
        56'b00000000000000000000000000000000101000010000001001111001,
        //tile 403
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 404
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 405
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 406
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 407
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 408
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 409
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 410
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 411
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 412
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 413
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 414
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 415
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 416
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 417
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 418
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 419
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 420
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 421
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 422
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 423
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 424
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 425
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 426
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 427
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 428
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 429
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 430
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 431
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 432
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 433
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 434
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 435
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 436
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 437
        56'b00000000000000000000000000000000000000101000001001110111,
        //tile 438
        56'b00000000000000000000000000000000000000001000101001111000,
        //tile 439
        56'b00000000000000000000000000000000101000010000001001111001,
        //tile 440
        56'b00000000000000000000000000000001000000101000001001111011,
        //tile 441
        56'b00000000000000000000000000000000000000001000101001111000,
        //tile 442
        56'b00000000000000000000000000000001000000101000001001111100,
        //tile 443
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 444
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 445
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 446
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 447
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 448
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 449
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 450
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 451
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 452
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 453
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 454
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 455
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 456
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 457
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 458
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 459
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 460
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 461
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 462
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 463
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 464
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 465
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 466
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 467
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 468
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 469
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 470
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 471
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 472
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 473
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 474
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 475
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 476
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 477
        56'b00000000000000000000000000000001000000101000001001111011,
        //tile 478
        56'b00000000000000000000000000000000000000001000101001111000,
        //tile 479
        56'b00000000000000000000000000000001000000101000001001111100,
        //tile 480
        56'b00000000000000000000000000000001000000101000001001111110,
        //tile 481
        56'b00000000000000000000000000000000000000001000101001111000,
        //tile 482
        56'b00000000000000000000000000000001000000101000001001111111,
        //tile 483
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 484
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 485
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 486
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 487
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 488
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 489
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 490
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 491
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 492
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 493
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 494
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 495
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 496
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 497
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 498
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 499
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 500
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 501
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 502
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 503
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 504
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 505
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 506
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 507
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 508
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 509
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 510
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 511
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 512
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 513
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 514
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 515
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 516
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 517
        56'b00000000000000000000000000000001000000101000001001111110,
        //tile 518
        56'b00000000000000000000000000000000000000001000101001111000,
        //tile 519
        56'b00000000000000000000000000000001000000101000001001111111,
        //tile 520
        56'b00000000000000000000000000000000000000101000001010000001,
        //tile 521
        56'b00000000000000000000000000000000000000101000001010000010,
        //tile 522
        56'b00000000000000000000000000000000000000101000001010000011,
        //tile 523
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 524
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 525
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 526
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 527
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 528
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 529
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 530
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 531
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 532
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 533
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 534
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 535
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 536
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 537
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 538
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 539
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 540
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 541
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 542
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 543
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 544
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 545
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 546
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 547
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 548
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 549
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 550
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 551
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 552
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 553
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 554
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 555
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 556
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 557
        56'b00000000000000000000000000000000000000101000001010000001,
        //tile 558
        56'b00000000000000000000000000000000000000101000001010000010,
        //tile 559
        56'b00000000000000000000000000000000000000101000001010000011,
        //tile 560
        56'b00000000000000000000000000001100000100010000001010000100,
        //tile 561
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 562
        56'b00000000000000000000000000001100000100001000010010000101,
        //tile 563
        56'b00000000000000000000000000000000000000101000001010000110,
        //tile 564
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 565
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 566
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 567
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 568
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 569
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 570
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 571
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 572
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 573
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 574
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 575
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 576
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 577
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 578
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 579
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 580
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 581
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 582
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 583
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 584
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 585
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 586
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 587
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 588
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 589
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 590
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 591
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 592
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 593
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 594
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 595
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 596
        56'b00000000000000000000000000000000000000101000001010001001,
        //tile 597
        56'b00000000000000000000000000001100000100010000001010000100,
        //tile 598
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 599
        56'b00000000000000000000000000001100000100001000010010000101,
        //tile 600
        56'b00000000000000000000000000001000001100000100010010001010,
        //tile 601
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 602
        56'b00000000000000000000000000001000001100000100010010001011,
        //tile 603
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 604
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 605
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 606
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 607
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 608
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 609
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 610
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 611
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 612
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 613
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 614
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 615
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 616
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 617
        56'b00000000000000000000000000001000001100000100010010001100,
        //tile 618
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 619
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 620
        56'b00000000000000000000000000001000001100000100010010001100,
        //tile 621
        56'b00000000000000000000000000001000001100000100010010001101,
        //tile 622
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 623
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 624
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 625
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 626
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 627
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 628
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 629
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 630
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 631
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 632
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 633
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 634
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 635
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 636
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 637
        56'b00000000000000000000000000001100000100010000001010001110,
        //tile 638
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 639
        56'b00000000000000000000000000001100000100010000001010001111,
        //tile 640
        56'b00000001111101000001101000001100010000001000000101011110,
        //tile 641
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 642
        56'b00000000000000000000000000001100010000001000000101011111,
        //tile 643
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 644
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 645
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 646
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 647
        56'b00000001111101000001101000001100010000001000000101011110,
        //tile 648
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 649
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 650
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 651
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 652
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 653
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 654
        56'b00000001111101000001101000001100010000001000000101011110,
        //tile 655
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 656
        56'b00111000001100111101001110000000010000001000000101001110,
        //tile 657
        56'b00000000110000001100101100001000110100000100010010010000,
        //tile 658
        56'b00000000001100110000101100001000000100010000110110010001,
        //tile 659
        56'b00000000110000001100101100001000110100000100010010010000,
        //tile 660
        56'b00000000001100110000101100001000000100010000110110010001,
        //tile 661
        56'b00111000001100111101001110000000010000001000000101001110,
        //tile 662
        56'b00000000111001001100111100001100010000001000000101001010,
        //tile 663
        56'b00000001111101000001101000001100010000001000000101011110,
        //tile 664
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 665
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 666
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 667
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 668
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 669
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 670
        56'b00000001111101000001101000001100010000001000000101100001,
        //tile 671
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 672
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 673
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 674
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 675
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 676
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 677
        56'b00000001111101000001101000001100010000001000000101100001,
        //tile 678
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 679
        56'b00000000000000000000000000001100010000001000000101011111,
        //tile 680
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 681
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 682
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 683
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 684
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 685
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 686
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 687
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 688
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 689
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 690
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 691
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 692
        56'b00000000000000000001100000001101100100001000000101100101,
        //tile 693
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 694
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 695
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 696
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 697
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 698
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 699
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 700
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 701
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 702
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 703
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 704
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 705
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 706
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 707
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 708
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 709
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 710
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 711
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 712
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 713
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 714
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 715
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 716
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 717
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 718
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 719
        56'b00000000000000000000000000001100010000001000000101100010,
        //tile 720
        56'b00000000000000000000000000001000000100001100010001100110,
        //tile 721
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 722
        56'b00000000000000000000000000001000000100001100010001100110,
        //tile 723
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 724
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 725
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 726
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 727
        56'b00000000000000000000000000001000000100001100010001100111,
        //tile 728
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 729
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 730
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 731
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 732
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 733
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 734
        56'b00000000000000000000000000001000000100001100010001100111,
        //tile 735
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 736
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 737
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 738
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 739
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 740
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 741
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 742
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 743
        56'b00000000000000000000000000001000000100001100010001100111,
        //tile 744
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 745
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 746
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 747
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 748
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 749
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 750
        56'b00000000000000000000000000001000000100001100010001101000,
        //tile 751
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 752
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 753
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 754
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 755
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 756
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 757
        56'b00000000000000000000000000001000000100001100010001101001,
        //tile 758
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 759
        56'b00000000000000000000000000001000000100001100010001101010,
        //tile 760
        56'b00000000000000000000000000001000001100000100010001101011,
        //tile 761
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 762
        56'b00000000000000000000000000001000000100001100010001101100,
        //tile 763
        56'b00000000000000000000000000000000101000001000010001101101,
        //tile 764
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 765
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 766
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 767
        56'b00000000000000000000000000000000101000010000001001110000,
        //tile 768
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 769
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 770
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 771
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 772
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 773
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 774
        56'b00000000000000000000000000000000101000010000001001110010,
        //tile 775
        56'b00000000000000010001011101011001010100101000001010010010,
        //tile 776
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 777
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 778
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 779
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 780
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 781
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 782
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 783
        56'b00000000000000000000000000000000101000010000001001110000,
        //tile 784
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 785
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 786
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 787
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 788
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 789
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 790
        56'b00000000000000000000000000000000101000010000001001110100,
        //tile 791
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 792
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 793
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 794
        56'b00000000000000000000000000000000000000101000001001101110,
        //tile 795
        56'b00000000000000000000000000000000000000101000001001101111,
        //tile 796
        56'b00000000000000000000000000000000000000101000001001110101,
        //tile 797
        56'b00000000000000000000000000001000001100000100010001110110,
        //tile 798
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 799
        56'b00000000000000000000000000001000000100001100010001101100,
        //tile 800
        56'b00000000000000000000000000000000000000101000001001110111,
        //tile 801
        56'b00000000000000000000000000000000000000001000101001111000,
        //tile 802
        56'b00000000000000000000000000000000101000010000001001111001,
        //tile 803
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 804
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 805
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 806
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 807
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 808
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 809
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 810
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 811
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 812
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 813
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 814
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 815
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 816
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 817
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 818
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 819
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 820
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 821
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 822
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 823
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 824
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 825
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 826
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 827
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 828
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 829
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 830
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 831
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 832
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 833
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 834
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 835
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 836
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 837
        56'b00000000000000000000000000000000000000101000001001110111,
        //tile 838
        56'b00000000000000000000000000000000000000001000101001111000,
        //tile 839
        56'b00000000000000000000000000000000101000010000001001111001,
        //tile 840
        56'b00000000000000000000000000000001000000101000001001111011,
        //tile 841
        56'b00000000000000000000000000000000000000001000101001111000,
        //tile 842
        56'b00000000000000000000000000000001000000101000001001111100,
        //tile 843
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 844
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 845
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 846
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 847
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 848
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 849
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 850
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 851
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 852
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 853
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 854
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 855
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 856
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 857
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 858
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 859
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 860
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 861
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 862
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 863
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 864
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 865
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 866
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 867
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 868
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 869
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 870
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 871
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 872
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 873
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 874
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 875
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 876
        56'b00000000000000000000000000000001000000101000001001111101,
        //tile 877
        56'b00000000000000000000000000000001000000101000001001111011,
        //tile 878
        56'b00000000000000000000000000000000000000001000101001111000,
        //tile 879
        56'b00000000000000000000000000000001000000101000001001111100,
        //tile 880
        56'b00000000000000000000000000000001000000101000001001111110,
        //tile 881
        56'b00000000000000000000000000000000000000001000101001111000,
        //tile 882
        56'b00000000000000000000000000000001000000101000001001111111,
        //tile 883
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 884
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 885
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 886
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 887
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 888
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 889
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 890
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 891
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 892
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 893
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 894
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 895
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 896
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 897
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 898
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 899
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 900
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 901
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 902
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 903
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 904
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 905
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 906
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 907
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 908
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 909
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 910
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 911
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 912
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 913
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 914
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 915
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 916
        56'b00000000000000000000000000000000101001000000001010000000,
        //tile 917
        56'b00000000000000000000000000000001000000101000001001111110,
        //tile 918
        56'b00000000000000000000000000000000000000001000101001111000,
        //tile 919
        56'b00000000000000000000000000000001000000101000001001111111,
        //tile 920
        56'b00000000000000000000000000000000000000101000001010000001,
        //tile 921
        56'b00000000000000000000000000000000000000101000001010000010,
        //tile 922
        56'b00000000000000000000000000000000000000101000001010000011,
        //tile 923
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 924
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 925
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 926
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 927
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 928
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 929
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 930
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 931
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 932
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 933
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 934
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 935
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 936
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 937
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 938
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 939
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 940
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 941
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 942
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 943
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 944
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 945
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 946
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 947
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 948
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 949
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 950
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 951
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 952
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 953
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 954
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 955
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 956
        56'b00000000000000000000000000000000000000101000001001111010,
        //tile 957
        56'b00000000000000000000000000000000000000101000001010000001,
        //tile 958
        56'b00000000000000000000000000000000000000101000001010000010,
        //tile 959
        56'b00000000000000000000000000000000000000101000001010000011,
        //tile 960
        56'b00000000000000000000000000001100000100010000001010000100,
        //tile 961
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 962
        56'b00000000000000000000000000001100000100001000010010000101,
        //tile 963
        56'b00000000000000000000000000000000000000101000001010000110,
        //tile 964
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 965
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 966
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 967
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 968
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 969
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 970
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 971
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 972
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 973
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 974
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 975
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 976
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 977
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 978
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 979
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 980
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 981
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 982
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 983
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 984
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 985
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 986
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 987
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 988
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 989
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 990
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 991
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 992
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 993
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 994
        56'b00000000000000000000000000000000000000101000001010000111,
        //tile 995
        56'b00000000000000000000000000000000000000101000001010001000,
        //tile 996
        56'b00000000000000000000000000000000000000101000001010001001,
        //tile 997
        56'b00000000000000000000000000001100000100010000001010000100,
        //tile 998
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 999
        56'b00000000000000000000000000001100000100001000010010000101,
        //tile 1000
        56'b00000000000000000000000000001000001100000100010010001010,
        //tile 1001
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1002
        56'b00000000000000000000000000001000001100000100010010010011,
        //tile 1003
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1004
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1005
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1006
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1007
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1008
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1009
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1010
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1011
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1012
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1013
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1014
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1015
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1016
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1017
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1018
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1019
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1020
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1021
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1022
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1023
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1024
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1025
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1026
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1027
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1028
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1029
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1030
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1031
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1032
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1033
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1034
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1035
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1036
        56'b00000000000000000000000000001000001100000100010000111000,
        //tile 1037
        56'b00000000000000000000000000001100000100010000001010001110,
        //tile 1038
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1039
        56'b00000000000000000000000000001100000100010000001010001110,
        //tile 1040
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1041
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1042
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1043
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1044
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1045
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1046
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1047
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1048
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1049
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1050
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1051
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1052
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1053
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1054
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1055
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1056
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1057
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1058
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1059
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1060
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1061
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1062
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1063
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1064
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1065
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1066
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1067
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1068
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1069
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1070
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1071
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1072
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1073
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1074
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1075
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1076
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1077
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1078
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1079
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1080
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1081
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1082
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1083
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1084
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1085
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1086
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1087
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1088
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1089
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1090
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1091
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1092
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1093
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1094
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1095
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1096
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1097
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1098
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1099
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1100
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1101
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1102
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1103
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1104
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1105
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1106
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1107
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1108
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1109
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1110
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1111
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1112
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1113
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1114
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1115
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1116
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1117
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1118
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1119
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1120
        56'b00000000000000000000100100100000011000010100011110010100,
        //tile 1121
        56'b00000000000000000000000000100100011000100000010110010101,
        //tile 1122
        56'b00000000000000000000000000100100011000100000010110010101,
        //tile 1123
        56'b00000000000000000000100100011000100000011100010110010110,
        //tile 1124
        56'b00000000000000000000000001011101011001010101010010010111,
        //tile 1125
        56'b00000000000000000000000001011101011001010101010010011000,
        //tile 1126
        56'b00000000000000000000000001011101011001010101010010011000,
        //tile 1127
        56'b00000000000000000000000001011101011001010101010010011000,
        //tile 1128
        56'b00000000000000000000000001011101011001010101010010011001,
        //tile 1129
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1130
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1131
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1132
        56'b10101010100110100000010010011100001100001000000110011010,
        //tile 1133
        56'b00000000000010011110100000010000001100001000000110011011,
        //tile 1134
        56'b00000000000010100000010010011100001100001000000110011100,
        //tile 1135
        56'b00000000000000010010100010011100001100001000000110011101,
        //tile 1136
        56'b00000000000000000000010010011100001100001000000110011110,
        //tile 1137
        56'b00000000000000000000010010011100001100001000000110011111,
        //tile 1138
        56'b00000000000010100000010010011100001100001000000110100000,
        //tile 1139
        56'b00000000000000000010100010011100001100001000000110100001,
        //tile 1140
        56'b00000010100110101010011100010000001100001000000110100010,
        //tile 1141
        56'b00000000000000000000010010011100001100001000000110100011,
        //tile 1142
        56'b00000000000000000010011100010000001100001000000110100100,
        //tile 1143
        56'b00000000000000000000000010011100001100001000000110100101,
        //tile 1144
        56'b00000000000000000000000010011100001100001000000110100110,
        //tile 1145
        56'b00000000000000000010100100010000001100001000000110100111,
        //tile 1146
        56'b00000000000000000010100100010000001100001000000110101000,
        //tile 1147
        56'b00000000000000000000100100100000011000010100011110010100,
        //tile 1148
        56'b00000000000000000000000000100100011000100000010110010101,
        //tile 1149
        56'b00000000000000000000000000100100011000100000010110010101,
        //tile 1150
        56'b00000000000000000000000000100100011000100000010110010101,
        //tile 1151
        56'b00000000000000000000100100011000100000011100010110010110,
        //tile 1152
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1153
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1154
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1155
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1156
        56'b00000000000000000000000000000000001100001000000100001000,
        //tile 1157
        56'b00000000000000000000000100101000001100010000001010101001,
        //tile 1158
        56'b00000000000000000000000100001100101000001000010010101010,
        //tile 1159
        56'b00000000000000000000000100001100101000001000010010101011,
        //tile 1160
        56'b00000000000000000000000000000000000000011000010110101100,
        //tile 1161
        56'b00000000000000000000000000001100000100010000001010101101,
        //tile 1162
        56'b00000000000000000000000000000000000000000000011010101110,
        //tile 1163
        56'b00000000000000000000000000000000000000010100011010101111,
        //tile 1164
        56'b00000000000000000000000001010001011101011001010110110000,
        //tile 1165
        56'b00000000000000000000000001010101011101011001010010110001,
        //tile 1166
        56'b00000000000000000000000001010101011101011001010010110001,
        //tile 1167
        56'b00000000000000000000000001010101011101011001010010110001,
        //tile 1168
        56'b00000000000000000000000001010101011101011001010010110010,
        //tile 1169
        56'b00000000000000000000000000001100000100010000001010110011,
        //tile 1170
        56'b00000000000000000000000000001100001000000100010010110100,
        //tile 1171
        56'b00000000000000000000000000001100000100001000010010110101,
        //tile 1172
        56'b00000000000000001110100010101110100110101000010010110110,
        //tile 1173
        56'b00000000000010101000010010101110100110011110100010110111,
        //tile 1174
        56'b00000000000000000010101010100100010010011110100010111000,
        //tile 1175
        56'b00000000000000000010101010100100010010100010011110111001,
        //tile 1176
        56'b00000010100110101010011110100000001000000100010010111010,
        //tile 1177
        56'b00000010101010100110011110100000010000001000000110111011,
        //tile 1178
        56'b00000000000000000010101010100110100010011100010010111100,
        //tile 1179
        56'b00000000000000000010100110101000010010100010011110111101,
        //tile 1180
        56'b00000000000000000010100010100100010010101010011110111110,
        //tile 1181
        56'b00000000000000000010100110100010101010011100010010111111,
        //tile 1182
        56'b00000000000000000010100010100110101010011100010011000000,
        //tile 1183
        56'b00000000000000000010101010100110100000010010011111000001,
        //tile 1184
        56'b00000000010010100000000100001010100110101010011111000010,
        //tile 1185
        56'b00000000000010011110100010101010100100010000000111000011,
        //tile 1186
        56'b00000000000000000000000000000000000000010010101011000100,
        //tile 1187
        56'b00000000000000000000000000000000000000011000010110101100,
        //tile 1188
        56'b00000000000000000000000000000000000000000000011010101110,
        //tile 1189
        56'b00000000000000000000000000000000000000000000011010101110,
        //tile 1190
        56'b00000000000000000000000000000000000000000000011010101110,
        //tile 1191
        56'b00000000000000000000000000000000000000010100011010101111,
        //tile 1192
        56'b00000000000000000000000001101101101001100101100011000101,
        //tile 1193
        56'b00000000000000000000000000000001101101101001100111000110,
        //tile 1194
        56'b00000000000000000000000000000001101101101001100111000110,
        //tile 1195
        56'b00000000000000000000000000000001101101101001100111000110,
        //tile 1196
        56'b00000000000000000000000001101101101001100001100111000111,
        //tile 1197
        56'b00000000000000000000000000101000001100000100010011001000,
        //tile 1198
        56'b00000000000000000000000000000000001100000100101011001001,
        //tile 1199
        56'b00000000000000000000000000010000001100000100101011001010
    
    };

    localparam bit [47:0] BITMAPS [3248] = '{


        // <--- FILE: MAP\CITY.PNG --->

        //tile 0, VRAM 56'b00000000000000000000000000010000001100001000000100000000
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011011011011011011011011011011011011011011011,
        //tile 1, VRAM 56'b00000000000000000000000000001100010000001000000100000001
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b000000000000000000000000000000000000000001000010,
        48'b001001001001001001001001001001001001001011000010,
        48'b000000000000000000000000000000000000000000000010,
        48'b001001001001001001001001001001001001001001001010,
        48'b011011011011011011011011011011011011011011011010,
        48'b010010010010010010010010010010010010010010010001,
        //tile 2, VRAM 56'b00000000000000000000100100100000011100011000010100000010
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001010000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000011011011011011011011011011011011011011011011,
        48'b000000000000000000000000000000000000000000000000,
        48'b000100100100100100100100100100100100100100100100,
        48'b000100100100100100100100100100100100100100100100,
        48'b000100100100100100100100100100100100100100100100,
        48'b000100100100100100100100100100100100100100100100,
        48'b000100100100100100100100100100100100100100100100,
        48'b000100100100100100100100100100100100100100100100,
        48'b010000000000000000000000000000000000000000000000,
        //tile 3, VRAM 56'b00000000000000000000000000100100100000010100011000000011
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b001001001001001001001001001001001001001001001001,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b001001001001001001001001001001001001001001001001,
        //tile 4, VRAM 56'b00000000000000000000100100100000011100010100011000000100
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b001001001001001001001001001001001001010000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b011011011011011011011011011011011011011011011001,
        48'b001001001001001001001001001001001001001001001001,
        48'b100100100100100100100100100100100100100100100001,
        48'b100100100100100100100100100100100100100100100001,
        48'b100100100100100100100100100100100100100100100001,
        48'b100100100100100100100100100100100100100100100001,
        48'b100100100100100100100100100100100100100100100001,
        48'b100100100100100100100100100100100100100100100001,
        48'b001001001001001001001001001001001001001001001010,
        //tile 5, VRAM 56'b00000000000000000000001000101000001100000100010000000101
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000010010010011010010010011010010010011010010010,
        48'b000010010010010010010010010010010010010010010010,
        48'b100100100000000100100000000100100000000100100000,
        //tile 6, VRAM 56'b00000000000000000000001000010000001100000100101000000110
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000010010010000010010010000010010010000010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b011100100011011100100011011100100011011100100011,
        //tile 7, VRAM 56'b00000000000000000000001000010000001100000100101000000111
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000010010010000010010010000010010010000010010011,
        48'b010010010010010010010010010010010010010010010011,
        48'b011100100011011100100011011100100011011100100100,
        //tile 8, VRAM 56'b00000000000000000000000000000000001100001000000100001000
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        //tile 9, VRAM 56'b00000000001000001100110100110000101100010000000100001001
        48'b000000001010011010011010011010011010011001100001,
        48'b000000001010011010011010011010011010011001100001,
        48'b000000001010011010011010011010011010011001100001,
        48'b101101001010011010011010011010011010011001100001,
        48'b000000001010011010011010011010011010011001100001,
        48'b000000001010011010011010011010011010011001100001,
        48'b000000001010011010011010011010011010011110001110,
        48'b101101001010011010011010011010011010011001000001,
        48'b000000001001001001001001001001001001001001001001,
        48'b000000001000000000000000000000000000000001110001,
        48'b000000110001001001001001001001001001001110110001,
        48'b101101001110110110110110110110110110110110110001,
        48'b000000001110001001001001001001001001001001110001,
        48'b000000001001110001001001001001001001001110001001,
        48'b000000001001110110001001001001001001110110001001,
        48'b101101001001001001001001001001001001001001001001,
        //tile 10, VRAM 56'b00000000000000000000000000001000001100000100010000001010
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000010010010010010010010010010010010010010010000,
        48'b000010011011011011011011011011011011011011010000,
        //tile 11, VRAM 56'b00000001001001000101000000111100101000010000111000001011
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000001010010001000000000,
        48'b000000011000000000000000001010100100010001001000,
        48'b000000000000000000001001001010100100010001011001,
        48'b011000000000000001011011001010001001010001000001,
        48'b000000000000000001000000000001000001001001001000,
        48'b000000000000000000001001001001001000000000000000,
        48'b000000000000101101000000000011000000000000000000,
        48'b000000000101110110101000000000000000000000000000,
        48'b011000101110100100110101000000000000000000000000,
        48'b000101110110100100110110101000000000000000000000,
        48'b000101110101110110101110101001001000000000000000,
        48'b000001101101110110101101011011011001000000000000,
        48'b001011011000101101001001000000001000000011000000,
        48'b001000000000001000000000001001000011011011000000,
        48'b000001001001000000000000000000000011011000000000,
        //tile 12, VRAM 56'b00000000000000000000000001001100111100111000010000001100
        48'b000001001001001001001010010010010010010010010010,
        48'b000001001001001001001001010010010010010010010010,
        48'b000001001001001001001001001010010010010010010011,
        48'b001000001001001001001001001010010010010010010011,
        48'b010001000011001001001011001001010010010010010010,
        48'b001001000001011011011001011001001010010010010010,
        48'b001001000001001001001001001011001010010010010010,
        48'b001001000001001001001001001001011001010010010010,
        48'b001001000001001001001001001001001011011011011010,
        48'b010001000001011001001001001001001001001001001011,
        48'b001001001000011001001001001001001001001001001001,
        48'b001001001001011011011011011001001001001001001001,
        48'b001001001001001000000011011011001001001001001001,
        48'b001001001001001010001000011011011011001001011001,
        48'b001001001001001001001001000011011011011011011001,
        48'b001001001001001001001001001000011011011011011011,
        //tile 13, VRAM 56'b00000000000000000000000000000001001100111000111100001101
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b010010010010001000000000000000000000000000000001,
        48'b000000000000010010010000000000000000000001010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000001000000000001,
        48'b000010010000000001000000000000001001001001001001,
        48'b010001001010010001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001010010010010,
        48'b010001001001001001001001001001001010001001001001,
        //tile 14, VRAM 56'b00000000000000000000000000010000111001001100111100001110
        48'b000000000000000000000001010010001010010010011010,
        48'b000000000000000000001010001001010010010010010011,
        48'b000000000000000010001010010010010010010010010011,
        48'b000000001000001001010010010010010010010010001011,
        48'b010001010001010010010010010010010010010001001011,
        48'b001010010010010010010010010010010010001001001011,
        48'b000010010010010010010010010010001001001001001011,
        48'b010010010010010010010010010001001001001001001011,
        48'b010010010010010010001010001001001001001001011010,
        48'b010010010010010010001001001001001001001011010010,
        48'b010010010010010010001001001001001001011010010010,
        48'b010010010010010001001001001011011011010010010010,
        48'b010001010010001001001001011010010010010010010010,
        48'b001010010001001001001011010010010010010000010010,
        48'b010010001001001001011010010010010000000000010010,
        48'b010001001001001011010010010010010000000010010010,
        //tile 15, VRAM 56'b00000000001000001100000100101100110000110100010000001111
        48'b000001000010011010011010011010011010011000100100,
        48'b000001000010011010011010011010011010011000100100,
        48'b000001000010011010011010011010011010011000100100,
        48'b000001000010011010011010011010011010011000101101,
        48'b000001000010011010011010011010011010011000100110,
        48'b000001000010011010011010011010011010011000100110,
        48'b110000110010011010011010011010011010011000100110,
        48'b000100000010011010011010011010011010011000101101,
        48'b000000000000000000000000000000000000000000100100,
        48'b000110000100100100100100100100100100100000100100,
        48'b000110110000000000000000000000000000000110100100,
        48'b000110110110110110110110110110110110110000101101,
        48'b000110000000000000000000000000000000110000100110,
        48'b000000110000000000000000000000000110000000100110,
        48'b000000110110000000000000000000110110000000100110,
        48'b000000000000000000000000000000000000000000101101,
        //tile 16, VRAM 56'b00000000000000000000000001011101011001010101010000010000
        48'b000001001000000001001000000001001000000001001000,
        48'b001010011001001010011001001010011001001010011001,
        48'b001001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b001010011000000010011000000010011000000010011000,
        48'b001010011000000010011000000010011000000010011000,
        48'b001001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b001010011000000010011000000010011000000010011000,
        48'b001010011000000010011000000010011000000010011000,
        48'b001001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b001010011000000010011000000010011000000010011000,
        48'b001010011000000010011000000010011000000010011000,
        48'b001001001000000001001000000001001000000001001000,
        48'b001001001001001001001001001001001001001001001001,
        //tile 17, VRAM 56'b00000000000000000000000001011101011001010101010000010001
        48'b000001001000000001001000000001001000000001001000,
        48'b001010011001001010011001001010011001001010011001,
        48'b000001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011000,
        48'b000010011000000010011000000010011000000010011000,
        48'b000001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011000,
        48'b000010011000000010011000000010011000000010011000,
        48'b000001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011000,
        48'b000010011000000010011000000010011000000010011000,
        48'b000001001000000001001000000001001000000001001000,
        48'b001001001001001001001001001001001001001001001001,
        //tile 18, VRAM 56'b00000000000000000000000001011101011001010101010000010010
        48'b000001001000000001001000000001001000000001001000,
        48'b001010011001001010011001001010011001001010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001001001001001001001001001001001001001001001001,
        //tile 19, VRAM 56'b00000000000000000000000001101101101001100101100000010011
        48'b000001001001001001001001001001001001001001001001,
        48'b001010010010010010010010010010010010010010010010,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001000001000001000001000001000001000001000001000,
        48'b000001001001001001001001001001001001001001001001,
        //tile 20, VRAM 56'b00000000000000000000000001100001101101101001100100010100
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000011000011000011000011000011000011000011000011,
        48'b000000000000000000000000000000000000000000000000,
        //tile 21, VRAM 56'b00000000000000000000000001101101101001100001100100010101
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001000001000001000001000001000001000001000000,
        48'b000000000000000000000000000000000000000000000001,
        //tile 22, VRAM 56'b00000000000000000000000000101000001100000100001000010110
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        //tile 23, VRAM 56'b00000000000000000000000000101000001100000100001000010111
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        //tile 24, VRAM 56'b00000000000000000000000000000001101101100001100100011000
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010001010010010010010010010010010010010010,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010010010010010010010010010001010010010010,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010010010001010010010010010010010010010010,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010010010010010010010010001010010010010010,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        //tile 25, VRAM 56'b00000000000000000000000000000001100101101101100000011001
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001000001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001000001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001000001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001000001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        //tile 26, VRAM 56'b00000000000000000000000000000001101101100101100000011010
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010000010010010010010010010010010010010001,
        48'b000000000000000000000000000000000000000000000001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010000010010010001,
        48'b000000000000000000000000000000000000000000000001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010000010010010010010010010010010001,
        48'b000000000000000000000000000000000000000000000001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010000010010010010001,
        48'b000000000000000000000000000000000000000000000001,
        48'b001001001001001001001001001001001001001001001001,
        //tile 27, VRAM 56'b00000000000000000000000001010101010001011101110000011011
        48'b000001001000001001001001001001001000001001001001,
        48'b000010010000010010010010010010010000010010010010,
        48'b000010010000010010010010010010010000010010010010,
        48'b000011011011011011011011011011011011011011011011,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011011,
        48'b000001001000001001001001001001001000001001001001,
        48'b000010010000010010010010010010010000010010010010,
        48'b000010010000010010010010010010010000010010010010,
        48'b000011011011011011011011011011011011011011011011,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011011,
        //tile 28, VRAM 56'b00000000000000000000000001010101010001110001011100011100
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010001010010010010010010010001010010010010,
        48'b010010010001010010010010010010010001010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010001010010010010010010010001010010010010,
        48'b010010010001010010010010010010010001010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011011,
        //tile 29, VRAM 56'b00000000000000000000000001010101010001110001011100011101
        48'b000000000001000000000000000000000001000000000001,
        48'b010010010001010010010010010010010001010010010001,
        48'b010010010001010010010010010010010001010010010001,
        48'b011011011011011011011011011011011011011011011001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011001,
        48'b000000000001000000000000000000000001000000000001,
        48'b010010010001010010010010010010010001010010010001,
        48'b010010010001010010010010010010010001010010010001,
        48'b011011011011011011011011011011011011011011011001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011001,
        //tile 30, VRAM 56'b00000000110000101100110100001100010000001000000100011110
        48'b000000000001000000000000000000000001000001010001,
        48'b000000000001000000000000000000000001000010000010,
        48'b000000000001000000000000000000000001000010010010,
        48'b011011011011011011011011011011011011011010100010,
        48'b000000001010010010010010010010010010010010100010,
        48'b000000010000000000000000000000000000000010100010,
        48'b000000010010010010010010010010010010010010100010,
        48'b011011010101110101110101110101110101110010100010,
        48'b000000010101110101110101110101110101110010100010,
        48'b000000010101110101110101110101110101110010100010,
        48'b000000010101110101110101110101110101110010100010,
        48'b011011010101110101110101110101110101110010100010,
        48'b000000010101110101110101110101110101110010100010,
        48'b000000010101110101110101110101110101110010100010,
        48'b000000010101110101110101110101110101110010100010,
        48'b011011010101110101110101110101110101110010100010,
        //tile 31, VRAM 56'b00000001000001001001000100111101001100010000111000011111
        48'b000000000000000000000000000000001001010010010010,
        48'b000000000000000000000000000000000000001001001001,
        48'b000000011000000000000000000000000000000000011000,
        48'b000000000000000000000000000000000000000000011011,
        48'b011000000000000011000000000000000000000000000011,
        48'b000000000000000011011011000000000000000000000000,
        48'b000000000000000000011011000000011000000000000000,
        48'b000000000000100100000000000011000000000000000000,
        48'b000000000100101101100000000000000000000000000000,
        48'b011000100101110110101100000000000000000000000000,
        48'b000100101101110110101101100000000000000000000000,
        48'b000100101100101101100101100001001000000000000000,
        48'b000001100100101101100100011011011001000000000000,
        48'b001011011000100100001001000000001000000011000000,
        48'b001000000000001000000000001001000011011011000000,
        48'b000001001001000000000000000000000011011000000000,
        //tile 32, VRAM 56'b00000000011100010101110000111100010000111001001100100000
        48'b000000000001001001001000000000000001001001001001,
        48'b010000000000000000001001001000001001001001000000,
        48'b010000000000000000000000000000000000000000000000,
        48'b001010000000010010000000000000000000000000010010,
        48'b011001010010100101010010000000000000000010001011,
        48'b001001001001100101101101010010010010010001001001,
        48'b001001001001100101101101101101101100001001001001,
        48'b001001001001100101101101101101101100001001001001,
        48'b001001001001100110101101101101110100001001001001,
        48'b011001100100110110110110110110110110100001001001,
        48'b100100101101110100100110100100110110110100001001,
        48'b100100100100100001100110100100100100101101100001,
        48'b001001001001001001100110100001001001100100001001,
        48'b001001001001001011100101100001001001001011001001,
        48'b001001001001001001100101100001001011011011001001,
        48'b001001001001001001001100001001001011011001001001,
        //tile 33, VRAM 56'b00000000000001000000111100101000111000010001001100100001
        48'b000000001001001010010010010010001001010010010010,
        48'b000001010010010010010010010001011011001010010010,
        48'b001010100010010010010010001011101101011001001010,
        48'b010010010010010010001001001011101101011001100001,
        48'b100010010010010001100100001011001001011001010001,
        48'b010010010010010001010010010001010001001001001010,
        48'b010010010010010010001001001001001010010010010010,
        48'b010010010010010010010010010100010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b100010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010100010010010010010010010100010010,
        48'b010010010010010010010010010010010100100100010010,
        48'b010010010010010010010010010010010100100010010010,
        //tile 34, VRAM 56'b00000000101100110000001100110100000100010000001000100010
        48'b000001000000010010010010010010010000010010010010,
        48'b001010001000010010010010010010010000010010010010,
        48'b001001001000010010010010010010010000010010010010,
        48'b001011001100100100100100100100100100100100100100,
        48'b001011001001001001001001001001001001001000010000,
        48'b001011001010010010010010010010010010010001010000,
        48'b001011001001001001001001001001001001001001010000,
        48'b001011001101110101110101110101110101110001100100,
        48'b001011001101110101110101110101110101110001010010,
        48'b001011001101110101110101110101110101110001010010,
        48'b001011001101110101110101110101110101110001010010,
        48'b001011001101110101110101110101110101110001100100,
        48'b001011001101110101110101110101110101110001010000,
        48'b001011001101110101110101110101110101110001010000,
        48'b001011001101110101110101110101110101110001010000,
        48'b001011001101110101110101110101110101110001100100,
        //tile 35, VRAM 56'b00000000000000000000000000010100011100100101110100100011
        48'b000001001000001001001001001001001000001001001001,
        48'b000010010000010010010010010010010000010010010010,
        48'b000010010000010010010010010010010000010010010010,
        48'b000011011011011011011011011011011011011011011011,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011011,
        48'b000001001000001001001001001001001000001001001001,
        48'b000010010000010010010010010010010000010010010010,
        48'b000010010000010010010010010010010000010010010010,
        48'b000011011011011011011011011011011011011011011011,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011011,
        //tile 36, VRAM 56'b00000000000000000000000000010100011101110100100100100100
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010001010010010010010010010001010010010010,
        48'b010010010001010010010010010010010001010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010001010010010010010010010001010010010010,
        48'b010010010001010010010010010010010001010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011011,
        //tile 37, VRAM 56'b00000000000000000000000000010100011101110100100100100101
        48'b000000000001000000000000000000000001000000000001,
        48'b010010010001010010010010010010010001010010010001,
        48'b010010010001010010010010010010010001010010010001,
        48'b011011011011011011011011011011011011011011011001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011001,
        48'b000000000001000000000000000000000001000000000001,
        48'b010010010001010010010010010010010001010010010001,
        48'b010010010001010010010010010010010001010010010001,
        48'b011011011011011011011011011011011011011011011001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010001010010010010010010010001,
        48'b010010010010010010010001010010010010010010010001,
        48'b011011011011011011011011011011011011011011011001,
        //tile 38, VRAM 56'b00000000000000000000101001111000001100000100001000100110
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001011011011011011011011011011011011001001,
        48'b000100100011011011011011011011011011001011100100,
        48'b000100100011011011011011011011011001001011100100,
        48'b000100100011011011011011011011001001011011100100,
        48'b000100100011011011011011011001001011011011100100,
        48'b000100100011011011011011001001011011011011100100,
        48'b000100100011011011011001001011011011011011100100,
        48'b000100100011011011001001011011011011001011100100,
        48'b000100100011011001001011011011011001011011100100,
        48'b000100100011001001011011011011001011011011100100,
        48'b000100100011001011011011011001011011011011100100,
        //tile 39, VRAM 56'b00000000000000000000101001111000001100000100001000100111
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001011011011011011011011011011011011001001,
        48'b100100100011011011011011011011011011001011100100,
        48'b100100100011011011011011011011011001001011100100,
        48'b100100100011011011011011011011001001011011100100,
        48'b100100100011011011011011011001001011011011100100,
        48'b100100100011011011011011001001011011011011100100,
        48'b100100100011011011011001001011011011011011100100,
        48'b100100100011011011001001011011011011001011100100,
        48'b100100100011011001001011011011011001011011100100,
        48'b100100100011001001011011011011001011011011100100,
        48'b100100100011001011011011011001011011011011100100,
        //tile 40, VRAM 56'b00000000000000000000000000101000001100000100001000101000
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        //tile 41, VRAM 56'b00000000000000000000000000101000001100000100001000101001
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 42, VRAM 56'b00000000000000000000101001111000001100000100001000101010
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001011011011011011011011011011011011001000,
        48'b100100100011011011011011011011011011001011100000,
        48'b100100100011011011011011011011011001001011100000,
        48'b100100100011011011011011011011001001011011100000,
        48'b100100100011011011011011011001001011011011100000,
        48'b100100100011011011011011001001011011011011100000,
        48'b100100100011011011011001001011011011011011100000,
        48'b100100100011011011001001011011011011001011100000,
        48'b100100100011011001001011011011011001011011100000,
        48'b100100100011001001011011011011001011011011100000,
        48'b100100100011001011011011011001011011011011100000,
        //tile 43, VRAM 56'b00000000001100010000111000000100111100101000001000101011
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001010010001001010010001001010010001001000,
        48'b000001001010010001001010010001001010010001001000,
        48'b000001001010010001001010010001001010010001001000,
        48'b000011011100100011011100100011011100100011011000,
        48'b000000000101101000000101101000000101101000000000,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101011101000000000000011011000000000011101011101,
        48'b101011101000000000011011000000000011000101011101,
        48'b101011101000000011011000000000011000000101011101,
        48'b101011101000011011000000000011000000000101011101,
        48'b101011000101101101101101101101101101101000011101,
        48'b101011000110110110110110110110110110110000011101,
        48'b101011011011011011011011011011011011011011011101,
        48'b000101101101101101101101101101101101101101101000,
        //tile 44, VRAM 56'b00000000000000000000101001111000001100000100001000101100
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001011011011011011011011011011011011001001000,
        48'b100100011011011011011011011011011001011100100000,
        48'b100100011011011011011011011011001001011100100000,
        48'b100100011011011011011011011001001011011100100000,
        48'b100100011011011011011011001001011011011100100000,
        48'b100100011011011011011001001011011011011100100000,
        48'b100100011011011011001001011011011011011100100000,
        48'b100100011011011001001011011011011001011100100000,
        48'b100100011011001001011011011011001011011100100000,
        48'b100100011001001011011011011001011011011100100000,
        48'b100100011011011011011011011011011011011100100000,
        //tile 45, VRAM 56'b00000000000000000000000000010000000100001001111000101101
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000001001001001001001001010010001001001000000,
        48'b000000001001001001001001010010001001001001000000,
        48'b000000011011011011011010010011011011011011000000,
        48'b000000011011011011010010011011011011011011000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000001001001001001001001010001001001001000000,
        48'b000000001001001001001001010001001001001001000000,
        48'b000000001001001001001010001001001001001001000000,
        48'b000000001001001001010001001001001001001001000000,
        48'b000000001001001010001001001001001001001001000000,
        48'b000000001001010001001001001001001001001001000000,
        48'b000000001010001001001001001001001001001001000000,
        48'b000000010001001001001001001011001001001011000000,
        //tile 46, VRAM 56'b00000000000000000000000000010000000100001001111000101110
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000001001001001001001001010010001001001000000,
        48'b000000001001001001001001010010001001001001000000,
        48'b000000011011011011011010010011011011011011000000,
        48'b000000011011011011010010011011011011011011000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000001001001001001001001010001001001001000000,
        48'b000000001001001001001001010001001001001001000000,
        48'b000000001001001001001010001001001001001001000000,
        48'b000000001001001001010001001001001001001001000000,
        48'b000000001001001010001001001001001001001001000000,
        48'b000000001001010001001001001001001001001001000000,
        48'b000000001010001001001001001001001001001001000000,
        48'b000000011001001001011001001001001001001001000000,
        //tile 47, VRAM 56'b00000000000000000000101001111000001100000100001000101111
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001011011011011011011011011011011011001001,
        48'b000100100011011011011011011011011011001011100100,
        48'b000100100011011011011011011011011001001011100100,
        48'b000100100011011011011011011011001001011011100100,
        48'b000100100011011011011011011001001011011011100100,
        48'b000100100011011011011011001001011011011011100100,
        48'b000100100011011011011001001011011011011011100100,
        48'b000100100011011011001001011011011011001011100100,
        48'b000100100011011001001011011011011001011011100100,
        48'b000100100011001001011011011011001011011011100100,
        48'b000100100011011011011011011011011011011011100100,
        //tile 48, VRAM 56'b00000000000000000000101001111000001100000100001000110000
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001011011011011011011011011011011011001000,
        48'b100100100011011011011011011011011011001011100000,
        48'b100100100011011011011011011011011001001011100000,
        48'b100100100011011011011011011011001001011011100000,
        48'b100100100011011011011011011001001011011011100000,
        48'b100100100011011011011011001001011011011011100000,
        48'b100100100011011011011001001011011011011011100000,
        48'b100100100011011011001001011011011011001011100000,
        48'b100100100011011001001011011011011001011011100000,
        48'b100100100011001001011011011011001011011011100000,
        48'b100100100011011011011011011011011011011011100000,
        //tile 49, VRAM 56'b00000000000000010000111000000100111100101000001000110001
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001010010001001010010001001010010001001010,
        48'b000001001010010001001010010001001010010001001010,
        48'b000001001010010001001010010001001010010001001010,
        48'b000011011100100011011100100011011100100011011100,
        48'b000000000101101000000101101000000101101000000101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101011101000011000000000000000000011000101011101,
        48'b101011101011000000000000000000011000000101011101,
        48'b101011101000000000000000000011000000000101011101,
        48'b101011101000000000000000011000000000000101011101,
        48'b101011101000000000000011000000000000000101011101,
        48'b101011101000000000011000000000000000000101011101,
        48'b101000101101101101101101101101101101101101000101,
        48'b101101011011011011011011011011011011011011101101,
        //tile 50, VRAM 56'b00000000000000010000000100111000101000111100001000110010
        48'b000000000000000000000000000000000000000000000000,
        48'b001010010001001010010001001010010001001010010000,
        48'b001010010001001010010001001010010001001010010000,
        48'b001010010001001010010001001010010001001010010000,
        48'b011100100011011100100011011100100011011100100000,
        48'b101000000101101000000101101000000101101000000000,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101100101000100000000000000000000100000101100101,
        48'b101100101100000000000000000000100000000101100101,
        48'b101100101000000000000000000100000000000101100101,
        48'b101100101000000000000000100000000000000101100101,
        48'b101100101000000000000100000000000000000101100101,
        48'b101100101000000000100000000000000000000101100101,
        48'b101000101101101101101101101101101101101101000101,
        48'b101101100100100100100100100100100100100100101101,
        //tile 51, VRAM 56'b00000000000000000001100001010001011001011101010100110011
        48'b000000000000000000000000000000000000000000000000,
        48'b000001010010010010010010010010010010010010001000,
        48'b000001000000000000000000000000000000000000001000,
        48'b000001000011011011011011011011011011011000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000000000000000000000000000000000000001000,
        48'b000001000000000000000000000000000000000000001000,
        48'b000001001001001001001001001001001001100100001000,
        //tile 52, VRAM 56'b00101100110000101000100001100001100100010000001000110100
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010001011011011011011011011011011011011011001010,
        48'b010001001001001001001001001001001001001001001010,
        48'b010001100100100101100101100101100100100100001010,
        48'b010001100100100100101100101100101100100100001010,
        48'b010001100100110101110101110101100100100100001010,
        48'b010001100110010010010010010010110110100100001010,
        48'b010001100110110110110110110110111100110100001010,
        48'b010001100100111110110110110111100111100100001010,
        48'b010001100111111111111111111111111100100100001010,
        48'b010001100111110110110110110110111100100100001010,
        48'b010001100100111111111111111111100100100100001010,
        48'b010001001001001001001001001001001001001001001010,
        48'b000001000000000000000000000000000000000000001000,
        48'b001001001001001001001001001001001001001001001001,
        //tile 53, VRAM 56'b00000000000000000000000001010101010001011101110000110101
        48'b000001001000001001001001001001001000001001001000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000011011011011011011011011011011011011011011000,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011000,
        48'b000001001000001001001001001001001000001001001000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000011011011011011011011011011011011011011011000,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011000,
        //tile 54, VRAM 56'b00000000000000000000000000001000001100000100101000110110
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011011011011011011011011011011011011011011011,
        //tile 55, VRAM 56'b00000000000000000000000000001000001100000100010000110111
        48'b000001001001001001001001001001001001001001001010,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000010001001001001001001001001001001001001001011,
        48'b011000001001001001001001001001001001001001001011,
        48'b011000010001001001001001001001001001001001001011,
        48'b011011000010010001001001001001001001001001001011,
        48'b011011011000000010010010010010010010010010010010,
        48'b011011011011011000000000000000000000000000000000,
        //tile 56, VRAM 56'b00000000000000000000000000001000001100000100010000111000
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        //tile 57, VRAM 56'b00000000000000000000000000001000010000000100001100111001
        48'b000001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001000010,
        48'b001001001001001001001001001001001001001001010011,
        48'b001001001001001001001001001001001001001000010011,
        48'b001001001001001001001001001001001000000010011011,
        48'b000000000000000000000000000000000010010011011011,
        48'b010010010010010010010010010010010011011011011011,
        //tile 58, VRAM 56'b01011001111100100101101000011101110100010000001000111010
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010001011010011011011011011011011010011011001010,
        48'b010001001001001001001001001001001001001001001010,
        48'b010001100100100100100101100100100100100100001010,
        48'b010001100100100100100011101101100100100100001010,
        48'b010001100100100100100110011011101101100100001010,
        48'b010001100100100100110110110110011011101100001010,
        48'b010001100100100100110111111110110110011101001010,
        48'b010001100100100110110111111110111110011100001010,
        48'b010001100100110111110110110110101011100100001010,
        48'b010001100100110110110110101011100100100100001010,
        48'b010001100110110110101011100100100100100100001010,
        48'b010001001001001001001001001001001001001001001010,
        48'b000001000000000000000000000000000000000000001000,
        48'b001001001001001001001001001001001001001001001001,
        //tile 59, VRAM 56'b01100001101101100100111000010000111100101000001000111011
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001010010001001010010001001010010001001010,
        48'b000001001010010001001010010001001010010001001010,
        48'b000001001010010001001010010001001010010001001010,
        48'b000011000100100011000100100011000100100011000100,
        48'b000000011011011000011011011000011011011000011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b101110101111111111111111111101110110110110110101,
        48'b101110101111111111111111111101110101101101110101,
        48'b101110101111111111111111111101110101111101110101,
        48'b101110101111111111111111111101110101111101110101,
        48'b101110101111111111111111111101110101101101110101,
        48'b101110101111111111111111111101110111111111110101,
        48'b101110101111111111111111111101110101101101110101,
        48'b101110101111111111111111111101110101111101110101,
        //tile 60, VRAM 56'b01100001101101100100010000111000101000111100001000111100
        48'b000000000000000000000000000000000000000000000000,
        48'b001010010001001010010001001010010001001010010000,
        48'b001010010001001010010001001010010001001010010000,
        48'b001010010001001010010001001010010001001010010000,
        48'b011100000011011100000011011100000011011100000000,
        48'b100000100100100000100100100000100100100000100000,
        48'b100100100100100100100100100100100100100100100100,
        48'b100100100100100100100100100100100100100100100100,
        48'b101110110110110110101111111111111111111101110101,
        48'b101110101101101110101111111111111111111101110101,
        48'b101110101111101110101111111111111111111101110101,
        48'b101110101111101110101111111111111111111101110101,
        48'b101110101101101110101111111111111111111101110101,
        48'b101110111111111110101111111111111111111101110101,
        48'b101110101101101110101111111111111111111101110101,
        48'b101110101111101110101111111111111111111101110101,
        //tile 61, VRAM 56'b00000001111000010000111000000100111100101000001000111101
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001010010001001010010001001010010001001010,
        48'b000001001010010001001010010001001010010001001010,
        48'b000001001010010001001010010001001010010001001010,
        48'b000011011100100011011100100011011100100011011100,
        48'b000000000101101000000101101000000101101000000101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b110110000000000000011000000000000000000000000000,
        48'b110110000000000011000000000000000000000000000011,
        48'b110110000000011000000000000000000000000000011011,
        48'b110110000011000000000000000000000000000011011000,
        48'b110110011101101101101101101101101101011011101101,
        48'b110110101101101101101101101101101011011101101101,
        48'b110110110110110110110110110110110110110110110110,
        48'b110110110110110110110110110110110110110110110110,
        //tile 62, VRAM 56'b00000001111000010000000100111000101000111100001000111110
        48'b000000000000000000000000000000000000000000000000,
        48'b001010010001001010010001001010010001001010010000,
        48'b001010010001001010010001001010010001001010010000,
        48'b001010010001001010010001001010010001001010010000,
        48'b011100100011011100100011011100100011011100100000,
        48'b101000000101101000000101101000000101101000000000,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b100100000000000000000000100000000000000000110110,
        48'b100000000000000000000100000000000000000000110110,
        48'b000000000000000000100000000000000000000000110110,
        48'b000000000000000100000000000000000000000000110110,
        48'b101101101101100101101101101101101101101101110110,
        48'b101101101100101101101101101101101101101101110110,
        48'b110110110110110110110110110110110110110110110110,
        48'b110110110110110110110110110110110110110110110110,
        //tile 63, VRAM 56'b00000000111001011101000001110100011100010000001000111111
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010001010011010010010010010010010011010010001011,
        48'b011001001001001001001001001001001001001001001011,
        48'b010001100100100100100100011011010010100100001011,
        48'b010001100100100100011010010010011011011100001011,
        48'b010001100100100010010011010011011011101110001011,
        48'b011001100100010011010010011011100101101110001011,
        48'b010001100010010010011011011100100011010010001011,
        48'b010001010010010011011101101110110010011011001011,
        48'b010001011011011100101101101011010010011100001011,
        48'b011001101110100100110011010010011011100100001011,
        48'b010001100110110010010010011011100100100100001011,
        48'b010001001001001001001001001001001001001001001011,
        48'b000001000000000000000000000000000000000000001000,
        48'b001001001001001001001001001001001001001001001001,
        //tile 64, VRAM 56'b01100001101101100100111000010000111100101000001001000000
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001010010001001010010001001010010001001000,
        48'b000001001010010001001010010001001010010001001000,
        48'b000001001010010001001010010001001010010001001000,
        48'b000011000100100011000100100011000100100011000000,
        48'b000000011011011000011011011000011011011000011000,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b101110101111111111111111111101110110110110110101,
        48'b101110101111111111111111111101110101101101110101,
        48'b101110101111111111111111111101110101111101110101,
        48'b101110101111111111111111111101110101111101110101,
        48'b101110101111111111111111111101110101101101110101,
        48'b101110101111111111111111111101110111111111110101,
        48'b101110101111111111111111111101110101101101110101,
        48'b101110101111111111111111111101110101111101110101,
        //tile 65, VRAM 56'b00000100101001000100110101100101100000010000001001000001
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010001010010010010010010010010010010010010001010,
        48'b011001001001001001001001001001001001001001001011,
        48'b010001100100100100100100101101101101100100001010,
        48'b010001100100100100100110101101101101101100001010,
        48'b010001100100100100100110110110101101101100001010,
        48'b011001100100100100110101110110110110111100001011,
        48'b010001100100100110110110110101111111101100001010,
        48'b010001100100100110101110111111111101101100001010,
        48'b010001100100110110111111111101101111101100001010,
        48'b011001100110111111111101101111101101100100001011,
        48'b010001100111111101101111101101100100100100001010,
        48'b010001001001001001001001001001001001001001001010,
        48'b000001000000000000000000000000000000000000001000,
        48'b001001001001001001001001001001001001001001001001,
        //tile 66, VRAM 56'b00000000000000000000000000000000001100001000000101000010
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        //tile 67, VRAM 56'b00000000000000000000000000000100010000001001111001000011
        48'b000000001001001001001001001010010010010010000000,
        48'b000000001001001001001001001000000000000000000000,
        48'b000000001001001001001001001001001001001011000000,
        48'b000000001001001001001001001001001001011011000000,
        48'b000000001001001001001001001001001011011001000000,
        48'b000000001001001001001001001001011011001001000000,
        48'b000000001001001001001001001011011001001001000000,
        48'b000000001001001001001001011011001001001011000000,
        48'b000000001001001001001011011001001001011001000000,
        48'b000000001001001001011011001001001011001001000000,
        48'b000000001001001011011001001001011001001001000000,
        48'b000000001001011011001001001011001001001001000000,
        48'b000000010011011010010010011010010010010010000000,
        48'b000000011011010010010011010010010010010010000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 68, VRAM 56'b00000000000000000000000000000100001000010001111001000100
        48'b000000001001001001001010010010010010010010000000,
        48'b000000000000000000000010010010010010010010000000,
        48'b000000010010010010010010010010010010010011000000,
        48'b000000010010010010010010010010010010011011000000,
        48'b000000010010010010010010010010010011011010000000,
        48'b000000010010010010010010010010011011010010000000,
        48'b000000010010010010010010010011011010010010000000,
        48'b000000010010010010010010011011010010010011000000,
        48'b000000010010010010010011011010010010011010000000,
        48'b000000010010010010011011010010010011010010000000,
        48'b000000010010010011011010010010011010010010000000,
        48'b000000010010011011010010010011010010010010000000,
        48'b000000001011011001001001011001001001001001000000,
        48'b000000011011001001001011001001001001001001000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 69, VRAM 56'b00000000000000000000000000000000001100000100001001000101
        48'b000001001001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010010010010010010010010010010010010010010,
        48'b000010010010010010010010010010010010010010010010,
        48'b000001001001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010010010010010010010010010010010010010010,
        48'b000010010010010010010010010010010010010010010010,
        48'b000001001001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010010010010010010010010010010010010010010,
        48'b000010010010010010010010010010010010010010010010,
        48'b000001001001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b000010010010010010010010010010010010010010010010,
        48'b000010010010010010010010010010010010010010010010,
        //tile 70, VRAM 56'b00000001101001010001000001100001011001011101010101000110
        48'b000001010010010010010010010010010011100100011000,
        48'b000001000000000000000000000000000011011011011000,
        48'b000001000101101101101101101101101011100100011000,
        48'b000001000001001001001001001001001011110110011000,
        48'b000001000001001001001001001001001001011011001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000001001001001001001001001001001000001000,
        48'b000001000000000000000000000000000000000000001000,
        48'b000001000000000000000000000000000000000000001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 71, VRAM 56'b00000000000000000000000000000001101101100001100101000111
        48'b000001001001001001001001001001001001001001001000,
        48'b000010010001010010010010010010010010010010010000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000010010010010010010010010010010001010010010000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000010010010010001010010010010010010010010010000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000010010010010010010010010010001010010010010000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 72, VRAM 56'b00000000110000001100101100110100000100010000001001001000
        48'b000001001001001001001001001001001001001001001001,
        48'b001010001011011011011011011011011011011011011011,
        48'b001001001000000000000000000000000000000000000000,
        48'b001000001100100100100100100100100100100100100100,
        48'b001000001100100100100100100100100100100100100100,
        48'b001001001000000000000000000000000000000000000000,
        48'b001101001110110110110110110110110110110110110110,
        48'b001101001100100100100100100100100100100100100100,
        48'b001101001110110110110110110110110110110110110110,
        48'b001001001000000000000000000000000000000000000000,
        48'b001000001100100100100100100100100100100100100100,
        48'b001001001001001001001001001001001001001001001001,
        48'b001000000001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b010010010010010010010000010010010010010010010000,
        48'b101101101101101101101101101101101101101101101101,
        //tile 73, VRAM 56'b00000000001100110000101100000100110100001000010001001001
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010000011000,
        48'b001001001001001001001001001001001001001000000000,
        48'b100100100100100100100100100100100100100000001000,
        48'b100100100100100100100100100100100100100000001000,
        48'b001001001001001001001001001001001001001000000000,
        48'b101101101101101101101101101101101101101000110000,
        48'b100100100100100100100100100100100100100000110000,
        48'b101101101101101101101101101101101101101000110000,
        48'b001001001001001001001001001001001001001000000000,
        48'b100100100100100100100100100100100100100000001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000000000001,
        48'b011011011011011011011001011011011011011011011001,
        48'b110110110110110110110110110110110110110110110110,
        //tile 74, VRAM 56'b00000000111001001100111100001100010000001000000101001010
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000010010010010000001000000000000,
        48'b011011011011011010100100100100010011011011011011,
        48'b000000000000010101110110110110101010000000000001,
        48'b000000000000001010101101101101010001000000000001,
        48'b000000000000010001010010010010001010000000000001,
        48'b011011011011010010010010010010010010011011011011,
        48'b000000000001010001011001001011001010000000000000,
        48'b000000000001010001011001001011001010000000000000,
        48'b000000000001010001011001001011001010000000000000,
        48'b011011011011011010001001001001010011011011011011,
        48'b000000000000000000010010010010000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b011011011011011011011011011011011011011011011011,
        //tile 75, VRAM 56'b00000000000000000000000000010100011100100101110101001011
        48'b000001001000001001001001001001001000001001001000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000011011011011011011011011011011011011011011000,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011000,
        48'b000001001000001001001001001001001000001001001000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000010010000010010010010010010010000010010010000,
        48'b000011011011011011011011011011011011011011011000,
        48'b000001001001001001001000001001001001001001001000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000010010010010010010000010010010010010010010000,
        48'b000011011011011011011011011011011011011011011000,
        //tile 76, VRAM 56'b00000000000000000000000000000001100001101101100101001100
        48'b000001000010010010010010010000001000010000001000,
        48'b000001000010010010010010010000001000000000001000,
        48'b000001000010010010010010010000001000010000001000,
        48'b000001000010010010010010010000001000000000001000,
        48'b000001000010010010010010010000001000000000001000,
        48'b000001000010010010010010010000001000000000001000,
        48'b000001000000000000000000000000001000000000001000,
        48'b000001000000000000000000000000001000010000001000,
        48'b000001001001001001001001001001001000000000001000,
        48'b000001000000000000000000000000001010010010001000,
        48'b000001000010010010010010010000001001001001001000,
        48'b000001000010010010010010010000001001001001001000,
        48'b000001000000000000000000000000001001001001001000,
        48'b000001000000000000000000000000001001001001001000,
        48'b000010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 77, VRAM 56'b00000000000000000000000000000001100001101101100101001101
        48'b000001000010000001000010010010010010010000001000,
        48'b000001000000000001000010010010010010010000001000,
        48'b000001000010000001000010010010010010010000001000,
        48'b000001000000000001000010010010010010010000001000,
        48'b000001000000000001000010010010010010010000001000,
        48'b000001000000000001000010010010010010010000001000,
        48'b000001000000000001000000000000000000000000001000,
        48'b000001000010000001000000000000000000000000001000,
        48'b000001000000000001001001001001001001001001001000,
        48'b000001010010010001000000000000000000000000001000,
        48'b000001001001001001000010010010010010010000001000,
        48'b000001001001001001000010010010010010010000001000,
        48'b000001001001001001000000000000000000000000001000,
        48'b000001001001001001000000000000000000000000001000,
        48'b000010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 78, VRAM 56'b00111000001100111101001110000000010000001000000101001110
        48'b000000000001000000010010010010000001000000000000,
        48'b000000000010010010011011011011010010010000000000,
        48'b000000010011011100101101101101100011011010000000,
        48'b110010011101101111100100100100111101101011010110,
        48'b010111100101101100101101101101100101101100111010,
        48'b010111101100100100111111111111100100100101111010,
        48'b000010101101101111100100100100111101101101010001,
        48'b010111100111111100101101101101100111111100111010,
        48'b010111101100100100111111111111100100100101111010,
        48'b000010101101101111100100100100111101101101010000,
        48'b000000010111111100111101101111100111111010000000,
        48'b110010111100100100111111111111100100100111010110,
        48'b010010111111111111100100100100111111111111010010,
        48'b010010010111111100111111111111100111111010010010,
        48'b010010010010010010111111111111010010010010010010,
        48'b110010010010010010010010010010010010010010010110,
        //tile 79, VRAM 56'b00000000000000000000000000001000001100000100010001001111
        48'b000001001001001001001001001001001001001001001010,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000010010010010010010010010010010010010010010010,
        48'b011000000000000000000000000000000000000000000000,
        //tile 80, VRAM 56'b00000000000000000000000000001000010000000100001101010000
        48'b000001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b000000000000000000000000000000000000000000000010,
        48'b010010010010010010010010010010010010010010010011,
        //tile 81, VRAM 56'b00000000000000000000000000001000001100000100010001010001
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001000,
        48'b000010010010010010010010010010010010010010010000,
        48'b011000000000000000000000000000000000000000000000,
        //tile 82, VRAM 56'b00000000000000000000000000001000001100000100010001010010
        48'b000001001001001001001001001001001001001001001010,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000010010010010010010010010010010010010010010011,
        48'b000010011011011011011011011011011011011011010011,
        //tile 83, VRAM 56'b00000000000000000000000000001000010000000100001101010011
        48'b000001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001010,
        48'b000000000000000000000000000000000000000000000010,
        48'b011000011011011011011011011011011011011011000010,
        //tile 84, VRAM 56'b00000010010010001110001010000100001100001000000101010100
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000011011011011011011011011011011011011011011011,
        48'b011100100100100100100101101101101101101101101101,
        48'b011100100011011011011011011011011011011011011100,
        48'b011100100011011011011011011011011011011011011100,
        48'b011100011101101101101101101101101101101101101100,
        48'b011100011101101101101101101101101101101101101100,
        48'b011100011101101101101101101101101101101101101100,
        48'b011101011101110110110110110110110110110110110100,
        48'b011101011101110110110110110110110110110110110100,
        48'b011101011101110110110110110110110110110110110100,
        48'b011101011101110110110110110110110110110110110100,
        //tile 85, VRAM 56'b00000000000010001010010110010010001110000100000101010101
        48'b000000000001001001001001001001001001001001001001,
        48'b000000001010010010010010010010010010010010010010,
        48'b000001010010011011011011011011011011011011011011,
        48'b001010100010011011011011011011011011011011011011,
        48'b001010100010011011011011011011011011011011011011,
        48'b010100100010011011011011011011011011011011011011,
        48'b100100100010011011011011011011011011011011011011,
        48'b100100100010011011011011011011011011011011011011,
        48'b100100100010011011011011011011011011011011011011,
        48'b100100100010011011011011011011011011011011011011,
        48'b100100100010011011011011011011011011011011011011,
        48'b100100100010011011011011011011011011011011011011,
        48'b100100100010011011011011011011011011011011011011,
        48'b100100100010010011011011011011011011011011011011,
        48'b100100100010010011011011011011011011011011011011,
        48'b100100101001001001001001001001001001001001001001,
        //tile 86, VRAM 56'b00000000000000000000000000000010010010001110000101010110
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        //tile 87, VRAM 56'b00000000000000000000000010010010001100000110000101010111
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 88, VRAM 56'b00111000111100001101000000101000010000001000000101011000
        48'b000000000001000000000000000000010010000000000000,
        48'b000000000001000000000000000010011011010000000000,
        48'b000000000001000000000000010011100100011010010000,
        48'b101101101101101101010010010011100100011010110010,
        48'b000000000000000010110110010011010010011010111010,
        48'b000000000000000010111111111010111010010010010001,
        48'b000000000000000000010010010010010000000000000001,
        48'b101101101101101101101101101101101101101101101101,
        48'b000000000001000010010000000000000001000000000000,
        48'b000000000001010011011010000000000001000000000000,
        48'b000000000010011100100011010010000001000000000000,
        48'b101010010010011100100011010110010101101101101101,
        48'b010110110010011010010011010111010000000000000001,
        48'b010111111111010111010010010010000000000000000001,
        48'b000010010010010010000001000000000000000000000001,
        48'b101101101101101101101101101101101101101101101101,
        //tile 89, VRAM 56'b00000000000000000000000000010000001100001000000101011001
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000011011000000000000001,
        48'b000000000000000000000001000011000000000000000001,
        48'b010010010010010010010010010011000011010010010010,
        //tile 90, VRAM 56'b00001000010000001100000110001010010010001110000101011010
        48'b000001000001010010010010010010010010010010010011,
        48'b000001000001010010010010010010010010010010010011,
        48'b000001000001010010010010010010010010010010010011,
        48'b000001000001001001001010010010010010010010010011,
        48'b000000000000000000000000000000000000000000000000,
        48'b000011011011011011011011011011011011011011011011,
        48'b000010010010010010010010010010010010010010010010,
        48'b000010010010010010010010010010010010010010010010,
        48'b000010010010010010010000000000000000000000000000,
        48'b000010010010010010010000000000000000000000000000,
        48'b100000000000000000000000011010010010010010010001,
        48'b101000010010010010000000000000000000000000000000,
        48'b100100000000000000000110110110100110100110100110,
        48'b100100110110110110110000000111111111111111111000,
        48'b100100110110110110110000000111111111111111111000,
        48'b101101101110110110110110110000000000000000000110,
        //tile 91, VRAM 56'b00000000010010011010010010000110001110001010010101011011
        48'b000001010010010010010010010010010010010010010010,
        48'b001010001011011010000000000000000000000000000010,
        48'b010100100011011010000000000000000000000000000010,
        48'b010100100011011010000000000000000000000000000010,
        48'b001011011011010010010010010010010010010010010011,
        48'b001100100011010001001001001001001001010010001011,
        48'b100100100011010001101101101101101101101101101011,
        48'b100100100011010001001001101101101101101101101011,
        48'b011100100011010001001001101101101101101101101011,
        48'b011100100011010001001001101101101101101101101011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011100100100100100100100100100100100100100100,
        48'b110011011011011011011011011011011011011011011011,
        48'b011110110110110110110110110110110110110110110110,
        48'b011110110110110110110110110110110110110110110110,
        48'b110110110110110110110110110110110110110110110110,
        //tile 92, VRAM 56'b00000000000000010000001010000110010010001010001101011100
        48'b000000000000000000000000000000000000000000000000,
        48'b001010010010010010010010010010010010010010010010,
        48'b001010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010011011,
        48'b010010010010010010010010010010010010010010011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b010010010010010010010010010010010010010010011011,
        48'b011011011011011011011011011011011011011011011100,
        48'b101101101101101101101101101101101101101101101011,
        48'b101101101101101101101101101101101101101101101011,
        48'b101101101101101101101101101101101101101101101101,
        //tile 93, VRAM 56'b00000000000000001000010000001110010010000110001101011101
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b010010010010010010010010010010010010010010010001,
        48'b001001001001001001001001001010010010010010010001,
        48'b001001001001001001001001001010010010010010010001,
        48'b000010010010010010010000001001001001001001001001,
        48'b001001001001001001001001001001010010010010001011,
        48'b100100011100011100011100100001001001001001100101,
        48'b001101101101101101101001001100100100100100100101,
        48'b001101101101101101101001001100100100100100100101,
        48'b100001001001001001001100100100100100100100011011,
        //tile 94, VRAM 56'b00000001111101000001101000001100010000001000000101011110
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000010010000000001000000000000,
        48'b000000000001000000010000000010000001000000000000,
        48'b011011011011011011010000000010011011011011011011,
        48'b000000000000000000010000000010000000000000000001,
        48'b000000000000000010000000000000010000000000000001,
        48'b000000000000000010000000000000010000000000000001,
        48'b011011011011011010011011011011010011011011011011,
        48'b000000000001000100010010010010100001000000000000,
        48'b000000000001000100101110110101100001000000000000,
        48'b000000000001000000100100100100000001000000000000,
        48'b011011011011011011010011011010011011011011011011,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b011011011011011011010011011010011011011011011011,
        //tile 95, VRAM 56'b00000000000000000000000000001100010000001000000101011111
        48'b000000000001000000000000000010000011010000000000,
        48'b000000000001000000000010010010010001010000000000,
        48'b000000000001000000010000000010010010000000000000,
        48'b011011011011011011010000000010010011010011011011,
        48'b000000000000000000010000000010010001010000000001,
        48'b000000000000000000010000000010010010000000000001,
        48'b000000000000000000010001001010010011010000000001,
        48'b011011011011011011010011011010010001010011011011,
        48'b000000000001000000001010010010010010000000000000,
        48'b000000000001000000010011011010010001000000000000,
        48'b000000000001000000010011011010010001000000000000,
        48'b011011011011011011010011011010011011011011011011,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b011011011011011011010011011010011011011011011011,
        //tile 96, VRAM 56'b00000000000000000000000000010000001100001000000101100000
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000011011000000000000000000001,
        48'b010010010010010010011010010011010010010010010010,
        48'b000000000001000000011010010011000001000000000000,
        48'b000000000001000000001011011001000001000000000000,
        48'b000000000001000000011001001011000001000000000000,
        48'b010010010010010010010011011010010010010010010010,
        48'b000000000000000000011000000011000000000000000001,
        48'b000000000000000000011011011011000000000000000001,
        48'b000000000000000000011001001011000000000000000001,
        48'b010010010010010010011001001011010010010010010010,
        //tile 97, VRAM 56'b00000001111101000001101000001100010000001000000101100001
        48'b000000000001000000000010010000000001000000000000,
        48'b000000000001000000010000000010000001000000000000,
        48'b000000000001000000010000000010000001000000000000,
        48'b011011011011011011010000000010011011011011011011,
        48'b000000000000000010000000000000010000000000000001,
        48'b000000000000000010000000000000010000000000000001,
        48'b000000000000000010011011011011010000000000000001,
        48'b011011011011011100010010010010100011011011011011,
        48'b000000000001000100101110110101100001000000000000,
        48'b000000000001000000100100100100000001000000000000,
        48'b000000000001000000010011011010000001000000000000,
        48'b011011011011011011010011011010011011011011011011,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b011011011011011011010011011010011011011011011011,
        //tile 98, VRAM 56'b00000000000000000000000000001100010000001000000101100010
        48'b000000000001000000010011011010000001000000000000,
        48'b000000000001000000010011011010000001000000000000,
        48'b000000000001000000010011011010000001000000000000,
        48'b011011011011011011010011011010011011011011011011,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b011011011011011011010011011010011011011011011011,
        48'b000000000001000000010011011010000001000000000000,
        48'b000000000001000000010011011010000001000000000000,
        48'b000000000001000000010011011010000001000000000000,
        48'b011011011011011011010011011010011011011011011011,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b000000000000000000010011011010000000000000000001,
        48'b011011011011011011010011011010011011011011011011,
        //tile 99, VRAM 56'b00000000000000000000000000010000001100001000000101100011
        48'b000000000001000000010011011010000001000000000000,
        48'b000000000001000000011000000011000001000000000000,
        48'b000000000001000000011011011011000001000000000000,
        48'b010010010010010010011001001011010010010010010010,
        48'b000000000000000000011001001011000000000000000001,
        48'b000000000000000000011001001011000000000000000001,
        48'b000000000000000000011001001011000000000000000001,
        48'b010010010010010010011001001011010010010010010010,
        48'b000000000001000000011001001011000001000000000000,
        48'b000000000001000000011001001011000001000000000000,
        48'b000000000001000000001011011001000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        //tile 100, VRAM 56'b00010001011100101001011000001101010100001000000101100100
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000010010000000001000000000000,
        48'b011011011011011011011010010011011011011011011011,
        48'b000000000000000000000010010000000000000000000001,
        48'b000000000000000000010100100010000000000000000001,
        48'b000000000000000000010101101010000000000000000001,
        48'b011011011011011011010101101010011011011011011011,
        48'b000000000001010010100100100100010010000000000000,
        48'b000000000010100010101100100101010100010000000000,
        48'b000000000010100010101101101101010100010000000000,
        48'b011011011010110110100101101100110110010011011011,
        48'b000000000111010010110110110110010010111000000001,
        48'b000000000000111111010010010010111111000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b011011011011011011011011011011011011011011011011,
        //tile 101, VRAM 56'b00000000000000000001100000001101100100001000000101100101
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000010010010010000001000000000000,
        48'b011011011011010010100100100100010010011011011011,
        48'b000000000010100100010010010010100100010000000001,
        48'b000000000010100010010100010100010100010000000001,
        48'b000000010100010010100010100010100010100010000001,
        48'b011011010100010100010100010100010010100010011011,
        48'b000000010100010010100010100010100010100010000000,
        48'b000000000010100010010100010100010100010000000000,
        48'b000000000010100100010010010010100100010000000000,
        48'b011011011011010010100100100100010010011011011011,
        48'b000000000000000000010010010010000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b011011011011011011011011011011011011011011011011,
        //tile 102, VRAM 56'b00000000000000000000000000001000000100001100010001100110
        48'b000000000000000000000001001000000000000000000000,
        48'b000010010010010010000001001000010010010010010001,
        48'b000010010010010010000001001000010010010010010011,
        48'b000010010010010010000001001000010010010010010011,
        48'b000010010010010010000001001000010010010010010011,
        48'b000010010010010010000001001000010010010010010000,
        48'b000010010010010000000001001000000010010010010000,
        48'b000010010010000001000001001000001000010010010000,
        48'b000010010000001001011001001011001001000010010000,
        48'b000010010010000011011011011011011000010010010000,
        48'b000010010010010000000000000000000010010010010000,
        48'b000010010010010010000000000000010010010010010000,
        48'b000010010010010010000000000000010010010010010000,
        48'b000010010010010010000000000000010010010010010000,
        48'b000001001001001001000000000000001001001001001000,
        48'b000001011011011011000000000000011011011011001000,
        //tile 103, VRAM 56'b00000000000000000000000000001000000100001100010001100111
        48'b000000000000000000000001001000000000000000000000,
        48'b010010010010010010000001001000010010010010010001,
        48'b010010010010010010000001001000010010010010010011,
        48'b010010010010010010000001001000010010010010010011,
        48'b010010010010010010000001001000010010010010010011,
        48'b010010010010010010000001001000010010010010010011,
        48'b010010010010010000000001001000000010010010010011,
        48'b010010010010000001000001001000001000010010010011,
        48'b010010010000001001011001001011001001000010010011,
        48'b010010010010000011011011011011011000010010010011,
        48'b010010010010010000000000000000000010010010010011,
        48'b010010010010010010000000000000010010010010010011,
        48'b010010010010010010000000000000010010010010010011,
        48'b010010010010010010000000000000010010010010010011,
        48'b001001001001001001000000000000001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        //tile 104, VRAM 56'b00000000000000000000000000001000000100001100010001101000
        48'b000000000000000000000001001000000000000000000000,
        48'b010010010010010010000001001000010010010010010001,
        48'b010010010010010010000001001000010010010010010011,
        48'b010010010010010010000001001000010010010010010011,
        48'b010010010010010010000001001000010010010010010011,
        48'b010010010010010000000001001000000010010010010011,
        48'b010010010010000001000001001000001000010010010011,
        48'b010010010000001001011001001011001001000010010011,
        48'b010010010010000011011011011011011000010010010011,
        48'b010010010010010000000000000000000010010010010011,
        48'b010010010010010010000000000000010010010010010011,
        48'b010010010010010010000000000000010010010010010011,
        48'b010010010010010010000000000000010010010010010011,
        48'b010010010010010010000000000000010010010010010011,
        48'b001001001001001001000000000000001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        //tile 105, VRAM 56'b00000000000000000000000000001000000100001100010001101001
        48'b000000000000000000000001001000000000000000000000,
        48'b010010010010010010000001001000010010010010010000,
        48'b010010010010010010000001001000010010010010010000,
        48'b010010010010010010000001001000010010010010010000,
        48'b010010010010010010000001001000010010010010010000,
        48'b010010010010010000000001001000000010010010010000,
        48'b010010010010000001000001001000001000010010010000,
        48'b010010010000001001011001001011001001000010010000,
        48'b010010010010000011011011011011011000010010010000,
        48'b010010010010010000000000000000000010010010010000,
        48'b010010010010010010000000000000010010010010010000,
        48'b010010010010010010000000000000010010010010010000,
        48'b010010010010010010000000000000010010010010010000,
        48'b010010010010010010000000000000010010010010010000,
        48'b001001001001001001000000000000001001001001001000,
        48'b000001011011011011000000000000011011011011001000,
        //tile 106, VRAM 56'b00000000000000000000000000001000000100001100010001101010
        48'b000000000000000000000001001000000000000000000000,
        48'b000010010010010010000001001000010010010010010001,
        48'b000010010010010010000001001000010010010010010011,
        48'b000010010010010010000001001000010010010010010011,
        48'b000010010010010010000001001000010010010010010011,
        48'b000010010010010010000001001000010010010010010011,
        48'b000010010010010000000001001000000010010010010011,
        48'b000010010010000001000001001000001000010010010011,
        48'b000010010000001001011001001011001001000010010011,
        48'b000010010010000011011011011011011000010010010011,
        48'b000010010010010000000000000000000010010010010011,
        48'b000010010010010010000000000000010010010010010011,
        48'b000010010010010010000000000000010010010010010011,
        48'b000010010010010010000000000000010010010010010011,
        48'b000001001001001001000000000000001001001001001001,
        48'b000001011011011011000000000000011011011011001000,
        //tile 107, VRAM 56'b00000000000000000000000000001000001100000100010001101011
        48'b000001001001001001000000000000001001001001001010,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000010001001001001000000000000001001001001001011,
        48'b011000001001001001001000000001001001001001001011,
        48'b011000010001001001001001001001001001001001001011,
        48'b011011000010010001001001001001001001001001001011,
        48'b011011011000000010010010010010010010010010010010,
        48'b011011011011011000000000000000000000000000000000,
        //tile 108, VRAM 56'b00000000000000000000000000001000000100001100010001101100
        48'b000001010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010010,
        48'b010010010010010010000000000000010010010010010001,
        48'b010010010010010010000000000000010010010010010000,
        48'b010010010010010010000000000000010010010010001000,
        48'b010010010010010010000000000000010010001001000011,
        48'b001001001001001001000000000000001001000000011011,
        48'b000000000000000000000000000000000000011011011011,
        //tile 109, VRAM 56'b00000000000000000000000000000000101000001000010001101101
        48'b000001001001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b000001010010010010010010010010010010010010010010,
        48'b000001010010010010010010010010010010010010010010,
        48'b000001010010001001001001001001001001001001001001,
        48'b000001010010001001001001001001001001001001001001,
        48'b000001010010001001001001001001001001001001001001,
        48'b000001010010001001001001001001001001001001001001,
        48'b000001010010001001001001001001001001001001001001,
        48'b000001010010001001001001001001001001001001001001,
        48'b000001010010001001001001001001001001001001001001,
        48'b001001010010001001001001001001001001001001001001,
        48'b001001010010010010001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001010010010010010010010010001001001001,
        //tile 110, VRAM 56'b00000000000000000000000000000000000000101000001001101110
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile 111, VRAM 56'b00000000000000000000000000000000000000101000001001101111
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001001001000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile 112, VRAM 56'b00000000000000000000000000000000101000010000001001110000
        48'b000000000000000000001001001001000000000000000000,
        48'b000000000000000000001001001001000000000000000000,
        48'b010010010010010010001001001001010010010010010010,
        48'b010010010010010010001001001001010010010010010010,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000000001001000000000000000000000,
        48'b010010010000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000010010010010010010010010000000000000,
        //tile 113, VRAM 56'b00000000000000000000000000000000000000101000001001110001
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile 114, VRAM 56'b00000000000000000000000000000000101000010000001001110010
        48'b000000000000000000001001001001000000000000000000,
        48'b000000000000000000001001001001000000000000000000,
        48'b010010010010010010001001001001010010010010010010,
        48'b010010010010010010001001001001010010010010010010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000000001001000000000000000000010,
        48'b000000000000000000000000000000000000000010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000010010010010010010010010000000000000,
        //tile 115, VRAM 56'b00000000000000000000000000000000101000010000001001110011
        48'b000000000000000000001001001001000000000000000000,
        48'b000000000000000000001001001001000000000000000000,
        48'b010010010010010010001001001001010010010010010010,
        48'b010010010010010010001001001001010010010010010010,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000001001001001000000000000000000,
        48'b010000000000000000000001001000000000000000000000,
        48'b010000000000000000000000000000000000000000000000,
        48'b010010010000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000010010010010010010010010000000000000,
        //tile 116, VRAM 56'b00000000000000000000000000000000101000010000001001110100
        48'b000000000000000000001001001001000000000000000000,
        48'b000000000000000000001001001001000000000000000000,
        48'b010010010010010010001001001001010010010010010010,
        48'b010010010010010010001001001001010010010010010010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000001001001001000000000000000010,
        48'b000000000000000000000001001000000000000000000010,
        48'b000000000000000000000000000000000000000000000010,
        48'b000000000000000000000000000000000000000010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000010010010010010010010010000000000000,
        //tile 117, VRAM 56'b00000000000000000000000000000000000000101000001001110101
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001000,
        48'b001001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile 118, VRAM 56'b00000000000000000000000000001000001100000100010001110110
        48'b000001001001001001000000000000001001001001001010,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000001001001001001000000000000001001001001001011,
        48'b000010001001001001001000000001001001001001001011,
        48'b011000001001001001001001001001001001001001001011,
        48'b011000010001001001001001001001001001001001001011,
        48'b011011000010010001001001001001001001001001001011,
        48'b011011011000000010010010010010010010010010010010,
        48'b011011011011011000000000000000000000000000000000,
        //tile 119, VRAM 56'b00000000000000000000000000000000000000101000001001110111
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile 120, VRAM 56'b00000000000000000000000000000000000000001000101001111000
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        //tile 121, VRAM 56'b00000000000000000000000000000000101000010000001001111001
        48'b000000000000000000001001001001000000000000000000,
        48'b000000000000010010001001001001010010000000000000,
        48'b000000000000010010001001001001010010000000000000,
        48'b000000000000010010001001001001000000000000000000,
        48'b000000000000010010001001001001000000000000000000,
        48'b000000000000010010000001001000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010000000000000000000000000000000,
        48'b000000000000010010010010010010010010000000000000,
        //tile 122, VRAM 56'b00000000000000000000000000000000000000101000001001111010
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile 123, VRAM 56'b00000000000000000000000000000001000000101000001001111011
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b010010010010010010010010010010001001000000000000,
        48'b010010010010010010010010010010001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        //tile 124, VRAM 56'b00000000000000000000000000000001000000101000001001111100
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001010010010010010010010010010010,
        48'b000000000000001001010010010010010010010010010010,
        48'b000000000000001001000000000000000000000000000000,
        //tile 125, VRAM 56'b00000000000000000000000000000001000000101000001001111101
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        //tile 126, VRAM 56'b00000000000000000000000000000001000000101000001001111110
        48'b000000000000000000000000000000001001000000000000,
        48'b010010010010010010010010010010001001000000000000,
        48'b010010010010010010010010010010001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile 127, VRAM 56'b00000000000000000000000000000001000000101000001001111111
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001010010010010010010010010010010,
        48'b000000000000001001010010010010010010010010010010,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile 128, VRAM 56'b00000000000000000000000000000000101001000000001010000000
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000010010010010010010010010000000000000,
        //tile 129, VRAM 56'b00000000000000000000000000000000000000101000001010000001
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000000000000000000000001001000000000000,
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 130, VRAM 56'b00000000000000000000000000000000000000101000001010000010
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        //tile 131, VRAM 56'b00000000000000000000000000000000000000101000001010000011
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 132, VRAM 56'b00000000000000000000000000001100000100010000001010000100
        48'b000000000000000001001001001001001001001001001001,
        48'b000000000001001010010010010010010010010010010011,
        48'b000000001010010010010010010010010010010010010000,
        48'b000001010010010010010010010010010010010010010000,
        48'b000001010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001011011011011011011011011011011011011011011000,
        48'b001011000000000000000000000000000000000000000011,
        //tile 133, VRAM 56'b00000000000000000000000000001100000100001000010010000101
        48'b000000000000000000000000000000000001001001001001,
        48'b010010010010010010010010010010010000000001001001,
        48'b010010010010010010010010010010010010010000001001,
        48'b010010010010010010010010010010010010010010000001,
        48'b010010010010010010010010010010010010010010000001,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011001001001001001001001001001001001001001011000,
        //tile 134, VRAM 56'b00000000000000000000000000000000000000101000001010000110
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000001001001001000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001000000000000000000000000000000000000000,
        48'b000001001001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 135, VRAM 56'b00000000000000000000000000000000000000101000001010000111
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000001001001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b000000000000000000000000000000000000000000000001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 136, VRAM 56'b00000000000000000000000000000000000000101000001010001000
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 137, VRAM 56'b00000000000000000000000000000000000000101000001010001001
        48'b000000000000001001001001001001001001000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000001001001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b000000000000000000000000000000000000000001001000,
        48'b001001001001001001001001001001001001001001001000,
        48'b001001001001001001001001001001001001001001001000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 138, VRAM 56'b00000000000000000000000000001000001100000100010010001010
        48'b000001001001001001001001001001001001001001001000,
        48'b010001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b011001001001001001001001001001001001001001001000,
        48'b010010010010010010010010010010010010010010010000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 139, VRAM 56'b00000000000000000000000000001000001100000100010010001011
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001010,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001000000001001001001011,
        48'b000010010010010010010010010000001010010010010010,
        48'b000000000000000000000000000000001000000000000000,
        //tile 140, VRAM 56'b00000000000000000000000000001000001100000100010010001100
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b010010010010010010010010010010010010010010010010,
        48'b011000000000000000000000000000000000000000000000,
        //tile 141, VRAM 56'b00000000000000000000000000001000001100000100010010001101
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001010,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b001001001001001001001001001001001001001001001011,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000011,
        //tile 142, VRAM 56'b00000000000000000000000000001100000100010000001010001110
        48'b000001001001001001001001001001001001001001001001,
        48'b001010010010010010010010010010010010010010010011,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001011011011011011011011011011011011011011011000,
        48'b001011000000000000000000000000000000000000000011,
        //tile 143, VRAM 56'b00000000000000000000000000001100000100010000001010001111
        48'b000001001001001001001001001001001001001001001001,
        48'b001010010010010010010010010010010010010010010011,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010010010010010010010000,
        48'b001010010010010010010010010001001010010010010000,
        48'b001011011011011011011011011001010011011011011000,
        48'b001011000000000000000000000001010001000000000011,
        //tile 144, VRAM 56'b00000000110000001100101100001000110100000100010010010000
        48'b000001000010010010010010010010010010010010010010,
        48'b000000000011011011011011011011011011011011011011,
        48'b000011000100100100100100100100100100100100100100,
        48'b000011000100100100100100100100100100100100100100,
        48'b000000000011011011011011011011011011011011011011,
        48'b000101000110110110110110110110110110110110110110,
        48'b000101000100100100100100100100100100100100100100,
        48'b000101000110110110110110110110110110110110110110,
        48'b000000000011011011011011011011011011011011011011,
        48'b000011000100100100100100100100100100100100100100,
        48'b000000000000000000000000000000000000000000000000,
        48'b000011011000000000000000000000000000000000000000,
        48'b011000000000000000000000000000000000000000000000,
        48'b001001001001001001001011001001001001001001001011,
        48'b001001001001001001001011001001001001001001001011,
        48'b101101101101101101101101101101101101101101101101,
        //tile 145, VRAM 56'b00000000001100110000101100001000000100010000110110010001
        48'b000000000000000000000000000000000000000001010001,
        48'b011011011011011011011011011011011011011001001001,
        48'b100100100100100100100100100100100100100001011001,
        48'b100100100100100100100100100100100100100001011001,
        48'b011011011011011011011011011011011011011001001001,
        48'b101101101101101101101101101101101101101001110001,
        48'b100100100100100100100100100100100100100001110001,
        48'b101101101101101101101101101101101101101001110001,
        48'b011011011011011011011011011011011011011001001001,
        48'b100100100100100100100100100100100100100001011001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001011011001,
        48'b001001001001001001001001001001001001001001001011,
        48'b010010010010010010010011010010010010010010010011,
        48'b010010010010010010010011010010010010010010010011,
        48'b110110110110110110110110110110110110110110110110,
        //tile 146, VRAM 56'b00000000000000010001011101011001010100101000001010010010
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001010010001001001001001001001,
        48'b001001001001001001001010010001001001001001001001,
        48'b001000000000000000000010010000000000000000000000,
        48'b001000000000000000010011011010000000000000000000,
        48'b001000000000000000010001001010000000000000000000,
        48'b001000000000000000010001001010000000000000000000,
        48'b001000000000010010011011011011010010000000000000,
        48'b001000000010011010001011011001010011010000000000,
        48'b001000000010011010001001001001010011010000000000,
        48'b001000000010100100011001001011100100010000000000,
        48'b001001001101010010100100100100010010101000000000,
        48'b000000000000101101010010010010101101000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000001001001001001001001001000000000000,
        //tile 147, VRAM 56'b00000000000000000000000000001000001100000100010010010011
        48'b000001001001001001001001001001001001001001001000,
        48'b000001001001001001001001001001001001001001001010,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000001001001001001001001001001001001001001001011,
        48'b000010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        //tile 148, VRAM 56'b00000000000000000000100100100000011000010100011110010100
        48'b000001001001001001001001001001001001001001001001,
        48'b001010011011011011011011011011011011011011011011,
        48'b001010010010010010010010010010010010010010010010,
        48'b001010010000001001001001001001001001001001001001,
        48'b001010010001100100100100100100100100100100100100,
        48'b001010010001100100100100100100100100100100100100,
        48'b001010010001100100100100100100100100100100100100,
        48'b001010010001100100100100100100100100100100100100,
        48'b001010010001100100100100100100100100100100100100,
        48'b001010010001100100100100100100100100100100100100,
        48'b001010010001001001001001001001001001001001001001,
        48'b001010010001010010010010010010010010010010010010,
        48'b001010010001010010010010010010010010010010010010,
        48'b001010010001010010010010010010010010010010010010,
        48'b001010010001010010010010010010010010010010010010,
        48'b001010010001010010010010010010010010010010010010,
        //tile 149, VRAM 56'b00000000000000000000000000100100011000100000010110010101
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b000000000000000000000000000000000000000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        //tile 150, VRAM 56'b00000000000000000000100100011000100000011100010110010110
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010000,
        48'b011011011011011011011011011011011011011011011000,
        48'b000000000000000000000000000000000000001011011000,
        48'b100100100100100100100100100100100100000011011000,
        48'b100100100100100100100100100100100100000011011000,
        48'b100100100100100100100100100100100100000011011000,
        48'b100100100100100100100100100100100100000011011000,
        48'b100100100100100100100100100100100100000011011000,
        48'b100100100100100100100100100100100100000011011000,
        48'b000000000000000000000000000000000000000011011000,
        48'b011011011011011011011011011011011011000011011000,
        48'b011011011011011011011011011011011011000011011000,
        48'b011011011011011011011011011011011011000011011000,
        48'b011011011011011011011011011011011011000011011000,
        48'b011011011011011011011011011011011011000011011000,
        //tile 151, VRAM 56'b00000000000000000000000001011101011001010101010010010111
        48'b000001001000000001001000000001001000000001001000,
        48'b001010011001001010011001001010011001001010011001,
        48'b001001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b001010011000000010011000000010011000000010011000,
        48'b001010011000000010011000000010011000000010011000,
        48'b001001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b001010011000000010011000000010011000000010011000,
        48'b001010011000000010011000000010011000000010011000,
        48'b001001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b001010011000000010011000000010011000000010011000,
        48'b001010011000000010011000000010011000000010011000,
        48'b001001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        //tile 152, VRAM 56'b00000000000000000000000001011101011001010101010010011000
        48'b000001001000000001001000000001001000000001001000,
        48'b001010011001001010011001001010011001001010011001,
        48'b000001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011000,
        48'b000010011000000010011000000010011000000010011000,
        48'b000001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011000,
        48'b000010011000000010011000000010011000000010011000,
        48'b000001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011000,
        48'b000010011000000010011000000010011000000010011000,
        48'b000001001000000001001000000001001000000001001000,
        48'b001000000001001000000001001000000001001000000001,
        //tile 153, VRAM 56'b00000000000000000000000001011101011001010101010010011001
        48'b000001001000000001001000000001001000000001001000,
        48'b001010011001001010011001001010011001001010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001000000001001000000001001000000001001000000001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000010011000000010011000000010011000000010011001,
        48'b000001001000000001001000000001001000000001001001,
        48'b001000000001001000000001001000000001001000000001,
        //tile 154, VRAM 56'b10101010100110100000010010011100001100001000000110011010
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000011000000001000000000000000000000001,
        48'b010010010011011011010010010010010010010010010010,
        48'b000000000001011000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000100100100000000000000,
        48'b010010010010010010010100100100100100100100100101,
        48'b000000000000000000100100100100110110110110100011,
        48'b000000000000100100100110110111110110100011101101,
        48'b000000000100100100110111111111110111011101101101,
        48'b100100100100111111110111111111110110110110101101,
        //tile 155, VRAM 56'b00000000000010011110100000010000001100001000000110011011
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000011011011011011000000000000000001000000000000,
        48'b011011011011011100100100100100100100010010010010,
        48'b100011011011101100100100100100100100100011011011,
        48'b100101101101101101101101100100100100100011011011,
        48'b100100101101101101101101101101100100100100011011,
        48'b100100100101101101101101101101101101101100011011,
        //tile 156, VRAM 56'b00000000000010100000010010011100001100001000000110011100
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010011010010010010010010010010010,
        48'b000000000001000011011011000000000001000000000000,
        48'b000000000001000000011000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b100000000000000000000001000000000000000000000001,
        48'b100100100100100100100100100000000000000000000001,
        48'b100100100100100100100100100100100100100000101101,
        48'b100100100100011101101101101101101100101101101101,
        //tile 157, VRAM 56'b00000000000000010010100010011100001100001000000110011101
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010011011011011011010010010010010010,
        48'b000000000000011011011011011011011000000000000001,
        48'b000000000000000011011011011011000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b100100100100100000000101101101101101101101101001,
        48'b100100100100100101101101101101101101101101101101,
        //tile 158, VRAM 56'b00000000000000000000010010011100001100001000000110011110
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000011,
        48'b000000000001000000000000000000000001000000011011,
        48'b000000000001000000000000000000000011011011011011,
        48'b010010010010010010010010010010011011011011011011,
        48'b000000000000000000000001000011011011011011011011,
        48'b000000000000000000000001000000011011011011011011,
        48'b000000000000000000000001000000000000011011011011,
        48'b100100100010010010010010010010010010010010010010,
        //tile 159, VRAM 56'b00000000000000000000010010011100001100001000000110011111
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011000001000000000000000000000001000000000000,
        48'b011011011001000000000000000000000001000000000000,
        48'b011011011011000000000000000000000001000000000000,
        48'b011011011010010010010010010010010010010010010100,
        48'b011011000000000000000001000100100100100100100100,
        48'b011000000000000000000100100100100100100100100100,
        48'b000000000000000000100100100100100100100100100100,
        48'b010010010010010100100100100100100100100100100100,
        //tile 160, VRAM 56'b00000000000010100000010010011100001100001000000110100000
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000011011011,
        48'b010010010010010010010010010010010011011011011011,
        48'b000000000001000000000000000011011011011011011011,
        48'b000000000001000000000000000011011011011011011011,
        48'b100100100100100100100000000011011011011011011011,
        48'b100100100100100100100100011011011011011011011011,
        48'b100100100100100100100011011011011011011011011011,
        48'b100100100100100100011011011011011011011011011011,
        48'b100100100100011011011011011101011011011011011011,
        48'b100100011011011011011101101101101011011011011011,
        //tile 161, VRAM 56'b00000000000000000010100010011100001100001000000110100001
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b011011000000000000000001000000000000000000000001,
        48'b011011011010010010010010010010010010010010010010,
        48'b011011011011011011000000000000000001000000000000,
        48'b011011011011011011011011011000000001011011011000,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011100011100011011011011011011011011011,
        48'b011011011100100100100100011011011011011011011011,
        //tile 162, VRAM 56'b00000010100110101010011100010000001100001000000110100010
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000011011011011000000000000000001000000000000,
        48'b100011011011011011011010010010010010010010010010,
        48'b100100011011011011011011000000000000000000000001,
        48'b100100011011101011011011011000000000000000011011,
        48'b100100100110101011100100100000000000000011011011,
        48'b100100110101101100100100100100100011011011011011,
        //tile 163, VRAM 56'b00000000000000000000010010011100001100001000000110100011
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000011000000000001000000000000000000000001,
        48'b000000011011011011011011000000000000000000000001,
        48'b010010011011011011011011011010010010010010010010,
        48'b000000000011011011011011000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000100100100100100100100100100100100100000001,
        48'b100100100100100100100100100100100100100100100100,
        48'b100100100100100100100100100100100100100100100100,
        48'b100100100100100100100100100100100100100100100100,
        //tile 164, VRAM 56'b00000000000000000010011100010000001100001000000110100100
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b011011000000000000000001000000000000000000000001,
        48'b011011011011011000100100100100100100100100100100,
        48'b011011011011100100100100100100100100100100100100,
        //tile 165, VRAM 56'b00000000000000000000000010011100001100001000000110100101
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b011011011000000000000001000000000000000000000001,
        48'b011011011011011011011011010010010010010010010010,
        //tile 166, VRAM 56'b00000000000000000000000010011100001100001000000110100110
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010011011011011011011011011011010010010010010010,
        //tile 167, VRAM 56'b00000000000000000010100100010000001100001000000110100111
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000011011011011011011011011000000001,
        48'b000000000000011011011011011011011011011011011011,
        48'b000000000011100100100100100100100100100011011011,
        48'b010010010011100100100100100100100100100100100100,
        //tile 168, VRAM 56'b00000000000000000010100100010000001100001000000110101000
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b000000000000000000000001000000000000000000000001,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b000000000001000000000000000000000001000000000000,
        48'b010010010010010010010010010010010010010010010010,
        48'b000000000000000000000001000000000000000000000001,
        48'b011011000000000000000001000000000000000000000001,
        48'b011011011011011011011011011011011000000000000001,
        48'b100011011011011011011011011011011011011011010010,
        //tile 169, VRAM 56'b00000000000000000000000100101000001100010000001010101001
        48'b000000000001001000000001001000000001001000000001,
        48'b001010010010011010010010011010010010011010010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        48'b001100010010011100010010011100010010011100010010,
        //tile 170, VRAM 56'b00000000000000000000000100001100101000001000010010101010
        48'b000001001000000001001000000001001000000001001000,
        48'b010011011011010011011011010011011011010011011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        48'b010100011011010100011011010100011011010100011011,
        //tile 171, VRAM 56'b00000000000000000000000100001100101000001000010010101011
        48'b000001001000000001001000000001001000000001001001,
        48'b010011011011010011011011010011011011010011011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        48'b010100011011010100011011010100011011010100011000,
        //tile 172, VRAM 56'b00000000000000000000000000000000000000011000010110101100
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        48'b000001001000001001001001001001001001001001001001,
        //tile 173, VRAM 56'b00000000000000000000000000001100000100010000001010101101
        48'b000001001001001001001001001001001001001001001000,
        48'b001010010001001000001001001001000001001010010001,
        48'b001010001000010001011011011011001000010001010001,
        48'b001001000010001011011011011011011001000010001001,
        48'b001000010000001011010010010010011001010000010001,
        48'b001000000010001010010010010010010001000010000001,
        48'b001000000000010001010010010010001000010000000001,
        48'b001001000011000010001001001001010000011000001001,
        48'b001000001000011000010000010000011000011001000001,
        48'b001011000001001000011000011000011001001000011001,
        48'b001011011000001001001001001001001001000011011001,
        48'b001011001001011011011011011011011011001001011001,
        48'b001001000000000000000000000000000000000000001001,
        48'b001011011011011011011011011011011011011011011001,
        48'b001011011011011011011011011011011011011011011001,
        48'b000001001001001001001001001001001001001001001000,
        //tile 174, VRAM 56'b00000000000000000000000000000000000000000000011010101110
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        //tile 175, VRAM 56'b00000000000000000000000000000000000000010100011010101111
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        48'b000000000000000000000000000000000000001000000001,
        //tile 176, VRAM 56'b00000000000000000000000001010001011101011001010110110000
        48'b000001010011011001010011011001010011011001010011,
        48'b000001010011011001010011011001010011011001010011,
        48'b000000000011011000000011011000000011011000000011,
        48'b000011011000000011011000000011011000000011011000,
        48'b000001010011011001010011011001010011011001010011,
        48'b000001010011011001010011011001010011011001010011,
        48'b000000000011011000000011011000000011011000000011,
        48'b000011011000000011011000000011011000000011011000,
        48'b000001010011011001010011011001010011011001010011,
        48'b000001010011011001010011011001010011011001010011,
        48'b000000000011011000000011011000000011011000000011,
        48'b000011011000000011011000000011011000000011011000,
        48'b000001010011011001010011011001010011011001010011,
        48'b000001010011011001010011011001010011011001010011,
        48'b000000000011011000000011011000000011011000000011,
        48'b000011011000000011011000000011011000000011011000,
        //tile 177, VRAM 56'b00000000000000000000000001010101011101011001010010110001
        48'b000001010000000001010000000001010000000001010000,
        48'b000001010000000001010000000001010000000001010000,
        48'b000011011000000011011000000011011000000011011000,
        48'b011000000011011000000011011000000011011000000011,
        48'b000001010000000001010000000001010000000001010000,
        48'b000001010000000001010000000001010000000001010000,
        48'b000011011000000011011000000011011000000011011000,
        48'b011000000011011000000011011000000011011000000011,
        48'b000001010000000001010000000001010000000001010000,
        48'b000001010000000001010000000001010000000001010000,
        48'b000011011000000011011000000011011000000011011000,
        48'b011000000011011000000011011000000011011000000011,
        48'b000001010000000001010000000001010000000001010000,
        48'b000001010000000001010000000001010000000001010000,
        48'b000011011000000011011000000011011000000011011000,
        48'b011000000011011000000011011000000011011000000011,
        //tile 178, VRAM 56'b00000000000000000000000001010101011101011001010010110010
        48'b000001010000000001010000000001010000000001010011,
        48'b000001010000000001010000000001010000000001010011,
        48'b000011011000000011011000000011011000000011011011,
        48'b011000000011011000000011011000000011011000000011,
        48'b000001010000000001010000000001010000000001010011,
        48'b000001010000000001010000000001010000000001010011,
        48'b000011011000000011011000000011011000000011011011,
        48'b011000000011011000000011011000000011011000000011,
        48'b000001010000000001010000000001010000000001010011,
        48'b000001010000000001010000000001010000000001010011,
        48'b000011011000000011011000000011011000000011011011,
        48'b011000000011011000000011011000000011011000000011,
        48'b000001010000000001010000000001010000000001010011,
        48'b000001010000000001010000000001010000000001010011,
        48'b000011011000000011011000000011011000000011011011,
        48'b011000000011011000000011011000000011011000000011,
        //tile 179, VRAM 56'b00000000000000000000000000001100000100010000001010110011
        48'b000001001001001001001001001001001001001001001001,
        48'b001010010010010010010010010010010010010010010010,
        48'b001010011000000000000000000000000000000000000000,
        48'b001010000011011011011011011011011011011011011011,
        48'b001010000000000000000000000000000000000000000000,
        48'b001010000011011011011011011011011011011011011011,
        48'b001010000011011011011011011011011011011011011011,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        48'b001010000010010010010010010010010010010010010010,
        //tile 180, VRAM 56'b00000000000000000000000000001100001000000100010010110100
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b010010010010010010010010010010010010010010010010,
        48'b011011011011011011011011011011011011011011011011,
        48'b011011011011011011011011011011011011011011011011,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        //tile 181, VRAM 56'b00000000000000000000000000001100000100001000010010110101
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010000,
        48'b001001001001001001001001001001001001001011010000,
        48'b011011011011011011011011011011011011011001010000,
        48'b001001001001001001001001001001001001001001010000,
        48'b011011011011011011011011011011011011011001010000,
        48'b011011011011011011011011011011011011011001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        48'b010010010010010010010010010010010010010001010000,
        //tile 182, VRAM 56'b00000000000000001110100010101110100110101000010010110110
        48'b000000001001001001001001001010010010010010010010,
        48'b000000001001001001001001001010010010010010010010,
        48'b000000001001001001001001001010001001010010011010,
        48'b000000001001001001001001001010010001001001001001,
        48'b000000001001001001001001001001010000000000001001,
        48'b000000001001001001001001001001010010000100100101,
        48'b000000001001001001001001001001010010011010100100,
        48'b000000001001001001001001001001001010010011010100,
        48'b000000001001001001001001001001001010010010011000,
        48'b000000001001001001001001001001001001010010010010,
        48'b000000001001001001001001001001001001010010010010,
        48'b000000001001001001001001001001001001001010010010,
        48'b000000001001001001001001001001001001001001010010,
        48'b000000001001001001001001001001001001001001001001,
        48'b000000001001001001001001001001001001001001001001,
        48'b000000001001001001001001001001001001001001001001,
        //tile 183, VRAM 56'b00000000000010101000010010101110100110011110100010110111
        48'b000000000000001001001001001001001000001001000000,
        48'b010000000000000000000000000000000000001000001001,
        48'b010010000000000000000000000000000000000001001001,
        48'b011010100000000000000000000000000000000000001001,
        48'b011010100000000000000000001001001000000000000000,
        48'b101010100000001101101000001000000000000000000001,
        48'b000100100000100100101101000000000000000000000000,
        48'b000000000000100100100000000000000000000000000000,
        48'b100000000000000000000000000000000100100100000000,
        48'b010010000000000000000000000100100100011000000000,
        48'b010010010100100100100100100010010010000000100100,
        48'b010010010010010010010010010010010010000000100101,
        48'b010010010010010010010010010010101101000000000101,
        48'b010010010010010010010010101101101101000000000000,
        48'b101101101101101101101101101101101100000000000000,
        48'b101101101101101101101101101101101000000000000000,
        //tile 184, VRAM 56'b00000000000000000010101010100100010010011110100010111000
        48'b000000000000000000000001001001000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001010010001001001001000001001001001001,
        48'b000001001001010010001001001000000000001001001001,
        48'b001000000000000000000011011011000000001001001001,
        48'b000000000000000010100100100100100000000001100011,
        48'b000000000000000010100100100100100100100010100100,
        48'b000001001000001010100100100100100100010010010100,
        48'b000001000001001010010100100100000000000000100100,
        48'b001000001001001001001100100100100000000000000000,
        48'b000001000001000001001001010100100000000010010000,
        48'b100100100000001000001001010000000000000010010000,
        48'b100100100100000000000000000000000000000000000000,
        48'b010100100100100010000000000000000000000000000000,
        48'b000000010100100010000000000000000000000000000011,
        48'b000000000000000000000000000000000000000000011011,
        //tile 185, VRAM 56'b00000000000000000010101010100100010010100010011110111001
        48'b000000000000000001010010010010010010010010010010,
        48'b000000000000000000010010010010010010010010010010,
        48'b000000000000000000000000010010010010010010010010,
        48'b000000000000000000000000000001000010010010010010,
        48'b000000000000000000000000000000001001001010010010,
        48'b011000000000000000000000000000000000001001001001,
        48'b100011010000000000000000000000000000000000000000,
        48'b100100000000000000000000000000010010010010010010,
        48'b100001000000000000000000010010010011011011011011,
        48'b001001001000000000000010010011011011011100100100,
        48'b001001000000000001001100100100100100100100100100,
        48'b001000001001001011011100100100100100100100100100,
        48'b001001000011100100100100100100100100100100100100,
        48'b001011100100100100100100100100100100100100100100,
        48'b011100100100100100100100100100100100100100100100,
        48'b100100100100100100100100100100100100100100100100,
        //tile 186, VRAM 56'b00000010100110101010011110100000001000000100010010111010
        48'b000000000000000001001001001001001010001001001001,
        48'b000000000000000000000001001001001010001001001001,
        48'b000000000000000000000000000001001011011011011011,
        48'b000000000000000000000011011011011011100011011011,
        48'b000000000000000011011011011011011011011011011011,
        48'b011011011011011011011011011000000011100100100000,
        48'b100100100100100100100100100000000100100011011101,
        48'b000100100100100100100100100100100011011101101101,
        48'b000000000000000000000000000000110110110101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        //tile 187, VRAM 56'b00000010101010100110011110100000010000001000000110111011
        48'b000000000001010010010010010010010010010010010010,
        48'b000000000010010010010010010010010010010010010010,
        48'b011011011011011010010010010010010010010010100100,
        48'b011011011011010010010101101101101101101101010010,
        48'b011010010010010101101101101101101101101101101101,
        48'b010010110110110110110110110110110110110110110110,
        48'b110110110110110110110110110110110110110110110110,
        48'b110110110110110110110110110110110110110110101101,
        48'b110110110110110110110110110110110110101101101101,
        48'b110110110110110110110110110110101101101101101101,
        48'b110110110110110110110110110101101101101101101101,
        48'b110110110110110110110110101101101101101101101010,
        48'b110110110110110110110110101101101101101101101010,
        48'b110110110110110110110110101101101101101101101101,
        48'b110110110110110110110110110110110110110110110110,
        48'b110110110110110110110110110110110110110110110110,
        //tile 188, VRAM 56'b00000000000000000010101010100110100010011100010010111100
        48'b000001001001001001010010010010010010001001001001,
        48'b000001001001001001010010010010010010010010010010,
        48'b001001001001001001010010010010010010010010010010,
        48'b000000000000000000000010010010010010010010010000,
        48'b011011011011011011011011010010010010010010010000,
        48'b100100100011011011011011011010001010010010010000,
        48'b011011011011011011010010010010001010010010010010,
        48'b011011011011011010010010010010010010010010010010,
        48'b011011011000000010010010010010010010010100100000,
        48'b011011011010010010010010010010010010010000100000,
        48'b011000010010010010010010010010010010010010010010,
        48'b000010010010010010010010010010010010010010010010,
        48'b000010010010010010010010010010010010010010010010,
        48'b000000000000000000000000000000000000000000000000,
        48'b100100100100100100100100100100100100100100100100,
        48'b100100100100100100100100100100100100100100100100,
        //tile 189, VRAM 56'b00000000000000000010100110101000010010100010011110111101
        48'b000001001001001001001001000000000000000000000000,
        48'b001001001001001001001001001000000000000000000000,
        48'b001001001001001001001001001001000000010000000000,
        48'b011011100100100001001001001001000000000000000000,
        48'b011011011011011010001001001000000000000000000000,
        48'b010010010010010001001001001000000000000000000001,
        48'b001001001001001001001001010001001001001010001010,
        48'b001001001001001001001001001001001001001010001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001010010010,
        48'b001001001001001001001001001001001001010100011100,
        48'b001001001001001001001001001001001010010100011011,
        48'b010010010010010010010010010010010010100100011011,
        48'b011011011011011011011011011011011011100100011011,
        48'b011011011011011011011011011011011011011011100011,
        //tile 190, VRAM 56'b00000000000000000010100010100100010010101010011110111110
        48'b000000001001001001001010010010010010010010010010,
        48'b000000010011001001001001001001011011011010010010,
        48'b000000010010011001001001001001001001011000000010,
        48'b000100000010010010010010001001001001000000000000,
        48'b100100100000000000000000000000000000000000000000,
        48'b100100100100000000000000000000000000000000000000,
        48'b100100100100000000000000000000000000000000000000,
        48'b100100100100000000000000000000000000100100100100,
        48'b100100100000100100100100100100100100100100100100,
        48'b100000000100010010010010010010010010010010010010,
        48'b010010010010010011011001001001001001001001001001,
        48'b011011011011011011011011001001001001001001001001,
        48'b001001001001001001001001011001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        //tile 191, VRAM 56'b00000000000000000010100110100010101010011100010010111111
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000000000000000000000000000,
        48'b000000000000000000000000001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001000000,
        48'b001001001001001001001001001001001000000000010010,
        48'b011011011011011011011011011011000000100100010010,
        48'b011011011011011011011011011011000100010010010010,
        48'b000000000000000000000011011000000100010010010010,
        48'b010010010010010100000000000000100010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        //tile 192, VRAM 56'b00000000000000000010100010100110101010011100010011000000
        48'b000000001001001001001001001001001001001001001001,
        48'b000001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b001001001001001001001001001001001001001001001001,
        48'b000000000000000001001001001001001001001001001001,
        48'b010010010010010000001001001001001001001001001001,
        48'b010010010010010010000001001001001001001001001001,
        48'b010010010010010010011000001001001001100100001001,
        48'b010010010010010010011000000000000000000100100100,
        48'b010010010010010010010011011011011010000000000100,
        48'b010010010010010010010010010010010010010010010000,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        //tile 193, VRAM 56'b00000000000000000010101010100110100000010010011111000001
        48'b000000000000000000000000000000001001001001001001,
        48'b000000000000000000000000000000000000001001000000,
        48'b000000000000000000000000000000000000000000000010,
        48'b000000000000000000000000000000000000000000000010,
        48'b000000000000000000000000000000000000000000000010,
        48'b000000000000000000000010010010010010010010010010,
        48'b000000000000000000010010010010010010010010010010,
        48'b000000000000000010010010010010010010010010010010,
        48'b000000000000010010010010000000000000000000010010,
        48'b010000000000010010010000000000000000000000000010,
        48'b010010010010010010000010000000000000000000010000,
        48'b001001010010010010010000010010000010000010000010,
        48'b011001001010010010010010010000010010010000010010,
        48'b100011001001001001001001010010010010010010010010,
        48'b100100011011011011001001001001001001010010010010,
        48'b100100100100100100011011011011011011001001001001,
        //tile 194, VRAM 56'b00000000010010100000000100001010100110101010011111000010
        48'b000000000000001010010010000000000011100100100100,
        48'b010000000001001001001001000000101000000000110110,
        48'b001001001001001110000000101101101101101101101101,
        48'b110110001001110110101101101101101101101101101101,
        48'b101110110001101101101101101101101101101101101101,
        48'b101101101101101101101101110101101101101000000101,
        48'b101101101101101101101101101101101000000000101000,
        48'b101101101101101101101101101101101000000000000101,
        48'b101101101101101101101101101101000000101000101101,
        48'b101101101101101101101101101000000101000101000101,
        48'b101101101101101101101110101101101000101000101101,
        48'b101101101101101101101101101101101101101101101110,
        48'b101101101101101101101101101101101101101101110110,
        48'b101101101101101101101101101101101101101101101101,
        48'b101101101101101101101101101101101101101101101101,
        48'b110101101101101101101101101101101101101101101101,
        //tile 195, VRAM 56'b00000000000010011110100010101010100100010000000111000011
        48'b000000000001010010010010010010010011011011011011,
        48'b001001001010010010011011011011011011011011011011,
        48'b001001001010010010011011011011011011011011011011,
        48'b100101001010010010010011011011011011011011011011,
        48'b100100001010010010010011011011011011011011011011,
        48'b100100001010010010010010011011011011011011011011,
        48'b100100001010010010010010010011011011011011011011,
        48'b100100001001010010010010010011011011011011011011,
        48'b100100100001001010010010010010011011011011011011,
        48'b100100100100001001001010010010010011011011011011,
        48'b100100100100100001001001010010010010011011011011,
        48'b100100100100100100100001001010010010010011011011,
        48'b100100100100100100100001010010010010010010011011,
        48'b100100100100001001001010010011011011011011011011,
        48'b100100001001010010010010011011011011011011011011,
        48'b001001010010010010011011011011011011011011011011,
        //tile 196, VRAM 56'b00000000000000000000000000000000000000010010101011000100
        48'b000000000000000000000000000000000000001001001001,
        48'b000000000000000000000000000000000000001001001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        48'b000000000000000000000000000000000000000000001001,
        //tile 197, VRAM 56'b00000000000000000000000001101101101001100101100011000101
        48'b000001001001001001001001001001001001001001001001,
        48'b001010010010010010010010010010010010010010010010,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        48'b001011011011011011011011011011011011011011011011,
        //tile 198, VRAM 56'b00000000000000000000000000000001101101101001100111000110
        48'b000000000000000000000000000000000000000000000000,
        48'b001001001001001001001001001001001001001001001001,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        48'b010010010010010010010010010010010010010010010010,
        //tile 199, VRAM 56'b00000000000000000000000001101101101001100001100111000111
        48'b000000000000000000000000000000000000000000000001,
        48'b010010010010010010010010010010010010010010010000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        48'b011011011011011011011011011011011011011011011000,
        //tile 200, VRAM 56'b00000000000000000000000000101000001100000100010011001000
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        48'b000001010010011001010010011001010010011001010010,
        //tile 201, VRAM 56'b00000000000000000000000000000000001100000100101011001001
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        48'b000001010010000001010010000001010010000001010010,
        //tile 202, VRAM 56'b00000000000000000000000000010000001100000100101011001010
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011,
        48'b000001010010000001010010000001010010000001010011
    
    };

    always_comb
    begin
        data      = DATA[Tile];
        bitmapIdx = 16 * data[7:0] + PixelY;
        bitmap    = BITMAPS[bitmapIdx];
        color     = bitmap[3*(15-PixelX) +: 3];
        Data      = data[6*color+8 +: 6];
    end

endmodule
