module text_pl_win_rom (
    input  logic PlayerTwo,
    input  logic [8:0] PixelX,
    input  logic [5:0] PixelY,
    output logic [5:0] Data
);

    logic [5:0] pixel;
    logic [47:0] data = 48'b00000000000000000000000111110000001000000101010;
    logic [980:0] bitmap;
    logic [2:0] color;

    localparam bit [980:0] BITMAPS [57] = '{


        // <--- FILE: ASSETS\TEXT\PL_WIN\WINNER.PNG --->

        //tile 0, VRAM 48'b000000000000000000000001111100000010000001010100
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001000000000000000000000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001000000000000000000000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001000000000000000000000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001000000000000000000000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001000000000000000000000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000001001001001001001001000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001000000000000000010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001000000000000000000000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000000000000000000000,
        981'b000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001000000000000000010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000001001001001001001,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000001001001001001001001001001001001001001001001001000000000000000000011011011011011011011011011011011011011011011011011011000000000000000011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011000000000000000000000000000000000001001001001001001,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000001001001001001001,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000001001001001001001,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000001001001001001001,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000001001001001001001,
        981'b000000000000000000010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000001001001001001001001001001001001000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000000001001001001001001,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001,
        981'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001,
        981'b001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000001001001001001001,
        981'b001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000001001001001001001,
        981'b001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000001001001001001001,
        981'b001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000001001001001001001,
        981'b001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000001001001001001001,
        981'b001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000000000001001001001001001
    
    };

    always_comb
    begin
        bitmap    = BITMAPS[0];
        color     = bitmap[3*(326-PixelX) +: 3];
        pixel     = data[6*color+0 +: 6];
        Data      = (0 < pixel && pixel < 6) ? pixel + PlayerTwo : pixel;
    end

endmodule
