module text_pl_anim_rom (
    input  logic PlayerTwo,
    input  logic [2:0] Tile,
    input  logic [6:0] PixelX,
    input  logic [7:0] PixelY,
    output logic [5:0] Data
);

    logic [5:0] pixel;
    logic [50:0] data;
    logic [11:0] bitmapIdx;
    logic [344:0] bitmap;
    logic [2:0] color;

    localparam bit [50:0] DATA [6] = '{


        // <--- FILE: ASSETS\TEXT\PL_ANIM\WIN.PNG --->

        //tile 0
        51'b111111101010010100000011000001110101110100000000000,
        //tile 1
        51'b111111101010010100000011000001110101110100000000001,
        //tile 2
        51'b111111101010010100000011000001110101110100000000010,
        //tile 3
        51'b111111101010010100000011000001110101110100000000011,
        //tile 4
        51'b111111101010010100000011000001110101110100000000100,
        //tile 5
        51'b111111101010010100000011000001110101110100000000101
    
    };

    localparam bit [344:0] BITMAPS [1350] = '{


        // <--- FILE: ASSETS\TEXT\PL_ANIM\WIN.PNG --->

        //tile 0, VRAM 51'b111111101010010100000011000001110101110100000000000
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        //tile 1, VRAM 51'b111111101010010100000011000001110101110100000000001
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        //tile 2, VRAM 51'b111111101010010100000011000001110101110100000000010
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110100100100100100100100100100100100011011011011011110110110110110110100100100100100011011011011011011011011011011011110110110110110110000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111000000000000000000000000000000000000000000000000,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000,
        //tile 3, VRAM 51'b111111101010010100000011000001110101110100000000011
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        //tile 4, VRAM 51'b111111101010010100000011000001110101110100000000100
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        //tile 5, VRAM 51'b111111101010010100000011000001110101110100000000101
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001010010010010010001001001001001001010010010010010001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001010010010010010001001001001001001010010010010010001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011100100100100100100001001001001001101101101101101101001001001001001011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100100100100100100010010010010010101101101101101101010010010010010100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000110110110110110011011011011011011011011011011011100100100100100100110110110110110011011011011011011100100100100100100100100100100100110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000111111111111111110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110111111111111111111111111111111111110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        345'b000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000
    
    };

    always_comb
    begin
        data      = DATA[Tile];
        bitmapIdx = 11'd225 * data[2:0] + PixelY;
        bitmap    = BITMAPS[bitmapIdx];
        color     = bitmap[3*(114-PixelX) +: 3];
        pixel     = data[6*color+3 +: 6];
        Data      = (0 < pixel && pixel < 6) ? pixel + PlayerTwo : pixel;
    end

endmodule
