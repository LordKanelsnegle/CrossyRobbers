module palette_rom (
    input logic [5:0] addr,
    output logic [23:0] data
);

    parameter bit [23:0] ROM [43] = '{
        24'b000000000000000000000000, //RGB(0,0,0)
        24'b101000111010011111000010, //RGB(163,167,194)
        24'b010000000100100101110011, //RGB(64,73,115)
        24'b011010000110111110011001, //RGB(104,111,153)
        24'b001011000011010101001101, //RGB(44,53,77)
        24'b010100100011001100111111, //RGB(82,51,63)
        24'b111111111010111001110000, //RGB(255,174,112)
        24'b100011110100110101010111, //RGB(143,77,87)
        24'b111111111100001010100001, //RGB(255,194,161)
        24'b101111010110101001100010, //RGB(189,106,98)
        24'b110111111110000011101000, //RGB(223,224,232)
        24'b010011000110100010000101, //RGB(76,104,133)
        24'b010011111010010010111000, //RGB(79,164,184)
        24'b100100101110100011000000, //RGB(146,232,192)
        24'b001110110111110101001111, //RGB(59,125,79)
        24'b011000111010101100111111, //RGB(99,171,63)
        24'b111100001011010101000001, //RGB(240,181,65)
        24'b110011000010111101111011, //RGB(204,47,123)
        24'b111001010110100010000011, //RGB(229,104,131)
        24'b001011110101011101010011, //RGB(47,87,83)
        24'b011110000001110101001111, //RGB(120,29,79)
        24'b010011110001110101001100, //RGB(79,29,76)
        24'b111001100100010100111001, //RGB(230,69,57)
        24'b101011010010111101000101, //RGB(173,47,69)
        24'b011111010011100000110011, //RGB(125,56,51)
        24'b001110110010000000100111, //RGB(59,32,39)
        24'b110011110111010100101011, //RGB(207,117,43)
        24'b101010110101000100110000, //RGB(171,81,48)
        24'b001010010001110100101011, //RGB(41,29,43)
        24'b001111010010100100110110, //RGB(61,41,54)
        24'b000101000001100000101110, //RGB(20,24,46)
        24'b111111111110111010000011, //RGB(255,238,131)
        24'b110010001101010001011101, //RGB(200,212,93)
        24'b000100010001000100010001, //RGB(17,17,17)
        24'b001111000011110000111100, //RGB(60,60,60)
        24'b000111100001111000011110, //RGB(30,30,30)
        24'b011001010111100101111101, //RGB(101,121,125)
        24'b000001100000011100001101, //RGB(6,7,13)
        24'b001001000001101100110011, //RGB(36,27,51)
        24'b000100100001010000101001, //RGB(18,20,41)
        24'b110010011101011111010011, //RGB(201,215,211)
        24'b100011111001110110011111, //RGB(143,157,159)
        24'b111011101110101011101010 //RGB(238,234,234)
    };

    assign data = ROM[addr];

endmodule