module money_rom (
    input  logic [1:0] Tile,
    input  logic [4:0] PixelX,
    input  logic [4:0] PixelY,
    output logic [5:0] Data
);

    logic [49:0] data;
    logic [6:0] bitmapIdx;
    logic [53:0] bitmap;
    logic [2:0] color;

    localparam bit [49:0] DATA [3] = '{


        // <--- FILE: ASSETS\MONEY\PALLETS.PNG --->

        //tile 0
        50'b00000000000000000001111111001111001000011100000000,
        //tile 1
        50'b01010001111111010001010111001111001000011100000001,
        //tile 2
        50'b11011001111111010111010011001111001000011100000010
    
    };

    localparam bit [53:0] BITMAPS [54] = '{


        // <--- FILE: ASSETS\MONEY\PALLETS.PNG --->

        //tile 0, VRAM 50'b00000000000000000001111111001111001000011100000000
        54'b000001010010010001010010010001010010010001010010010000,
        54'b000011010010010011010010010011010010010011010010010011,
        54'b001011010010010011010010010011010010010011010010010011,
        54'b001011010010010011010010010011010010010011010010010011,
        54'b001100010010010100010010010100010010010100010010010100,
        54'b000011010010010011010010010011010010010011010010010011,
        54'b001011010010010011010010010011010010010011010010010011,
        54'b001011010010010011010010010011010010010011010010010011,
        54'b001100010010010100010010010100010010010100010010010100,
        54'b000011010010010011010010010011010010010011010010010011,
        54'b001011010010010011010010010011010010010011010010010011,
        54'b001011010010010011010010010011010010010011010010010011,
        54'b001100010010010100010010010100010010010100010010010100,
        54'b000011010010010011010010010011010010010011010010010011,
        54'b001011010010010011010010010011010010010011010010010011,
        54'b001011010010010011010010010011010010010011010010010011,
        54'b001100011011011100011011011100011011011100011011011100,
        54'b000001001001000001001001000001001001000001001001000000,
        //tile 1, VRAM 50'b01010001111111010001010111001111001000011100000001
        54'b000001010010010001010010010001010010010001010010010000,
        54'b000011010010010011100100100011100100100011010010010011,
        54'b001011010010100100100100100100100100100100100010010011,
        54'b001011010010100100101101101100101101101100100010010011,
        54'b001110010010101101100100100101100100100101101010010110,
        54'b000011010010100100100100100100100100100100100010010011,
        54'b001011010010100100111111111100111111111100100010010011,
        54'b001011010010111111111010111111111010111111111010010011,
        54'b001110010010010110100100100110100100100110010010010110,
        54'b000011010010100100100100100100100100100100100010010011,
        54'b001011010010100100101101101100101101101100100010010011,
        54'b001011010010101101100100100101100100100101101010010011,
        54'b001110010010100100100100100100100100100100100010010110,
        54'b000011010010100100111111111100111111111100100010010011,
        54'b001011010010111111111010111111111010111111111010010011,
        54'b001011010010010011010010010011010010010011010010010011,
        54'b001110011011011110011011011110011011011110011011011110,
        54'b000001001001000001001001000001001001000001001001000000,
        //tile 2, VRAM 50'b11011001111111010111010011001111001000011100000010
        54'b000001010010010001010010010001010010010001010010010000,
        54'b000011010010010011100100010100100010100100010010010011,
        54'b001011010010101101100100101100100101100100101010010011,
        54'b001011010010101101100100101100100101100100101010010011,
        54'b001001010010101101100100101100100101100100101010010110,
        54'b000011010010101101100100101100100101100100101010010011,
        54'b001011010010101101111111101111111101111111101010010011,
        54'b001011010010111111010111111011111111010111111010010011,
        54'b001001010010010100100010100100010100100110010010010110,
        54'b000011010010101100100101100100101100100101101010010011,
        54'b001011010010101100100101100100101100100101101010010011,
        54'b001011010010101100100101100100101100100101101010010011,
        54'b001001010010101100100101100100101100100101101010010110,
        54'b000011010010101111111101111111101111111101101010010011,
        54'b001011010010111111010111111011111111010111111010010011,
        54'b001011010010010011010010010011010010010011010010010011,
        54'b001001011011011001011011011001011011011001011011011110,
        54'b000001001001000001001001000001001001000001001001000000
    
    };

    always_comb
    begin
        data      = DATA[Tile];
        bitmapIdx = 6'd18 * data[1:0] + PixelY;
        bitmap    = BITMAPS[bitmapIdx];
        color     = bitmap[3*(17-PixelX) +: 3];
        Data      = data[6*color+2 +: 6];
    end

endmodule
