module player_rom (
    input  logic PlayerTwo,
    input  logic [6:0] Tile,
    input  logic [4:0] PixelX,
    input  logic [4:0] PixelY,
    output logic [5:0] Data
);

    logic [5:0] pixel;
    logic [53:0] data;
    logic [10:0] bitmapIdx;
    logic [95:0] bitmap;
    logic [2:0] color;

    localparam bit [53:0] DATA [128] = '{


        // <--- FILE: ASSETS\PLAYER\1-IDLE.PNG --->

        //tile 0
        54'b101000111101111100000101101010000001000011000000000000,
        //tile 1
        54'b101000111100111101000101101010000001000011000000000001,
        //tile 2
        54'b101000111101000101101010111100000001000011000000000010,
        //tile 3
        54'b101000000101101010111101111100000001000011000000000011,
        //tile 4
        54'b101000111101111100000101101010000001000011000000000000,
        //tile 5
        54'b101000111100111101000101101010000001000011000000000001,
        //tile 6
        54'b101000111101000101101010111100000001000011000000000010,
        //tile 7
        54'b101000000101101010111101111100000001000011000000000011,
        //tile 8
        54'b101000111101111100000101101010000001000011000000000100,
        //tile 9
        54'b101000111100111101000101101010000001000011000000000101,
        //tile 10
        54'b101000111101111100000101101010000001000011000000000110,
        //tile 11
        54'b101000111101000101101010111100000001000011000000000111,
        //tile 12
        54'b101000111101111100000101101010000001000011000000001000,
        //tile 13
        54'b101000111100111101000101101010000001000011000000001001,
        //tile 14
        54'b101000111101111100000101101010000001000011000000001010,
        //tile 15
        54'b101000111101000101101010111100000001000011000000001011,
        //tile 16
        54'b101000111101111100000101101010000001000011000000001000,
        //tile 17
        54'b101000111100111101000101101010000001000011000000001001,
        //tile 18
        54'b101000111101111100000101101010000001000011000000001010,
        //tile 19
        54'b101000111101000101101010111100000001000011000000001011,
        //tile 20
        54'b101000111101111100000101101010000001000011000000000100,
        //tile 21
        54'b101000111100111101000101101010000001000011000000000101,
        //tile 22
        54'b101000111101111100000101101010000001000011000000000110,
        //tile 23
        54'b101000111101000101101010111100000001000011000000000111,
        //tile 24
        54'b101000111101111100000101101010000001000011000000000000,
        //tile 25
        54'b101000111100111101000101101010000001000011000000000001,
        //tile 26
        54'b101000111101000101101010111100000001000011000000000010,
        //tile 27
        54'b101000000101101010111101111100000001000011000000000011,
        //tile 28
        54'b101000111101111100000101101010000001000011000000000000,
        //tile 29
        54'b101000111100111101000101101010000001000011000000000001,
        //tile 30
        54'b101000111101000101101010111100000001000011000000000010,
        //tile 31
        54'b101000000101101010111101111100000001000011000000000011,

        // <--- FILE: ASSETS\PLAYER\2-WALK.PNG --->

        //tile 0
        54'b101000111101111100000101101010000001000011000000001100,
        //tile 1
        54'b101000111100111101000101101010000001000011000000001101,
        //tile 2
        54'b101000111101000101101010111100000001000011000000001110,
        //tile 3
        54'b101000000101101010111101111100000001000011000000001111,
        //tile 4
        54'b101000111101111100000101101010000001000011000000000000,
        //tile 5
        54'b101000111100111101000101101010000001000011000000000001,
        //tile 6
        54'b101000111101000101101010111100000001000011000000000010,
        //tile 7
        54'b101000000101101010111101111100000001000011000000000011,
        //tile 8
        54'b101000111101111100000101101010000001000011000000010000,
        //tile 9
        54'b101000111100111101000101101010000001000011000000010001,
        //tile 10
        54'b101000111101000101101010111100000001000011000000010010,
        //tile 11
        54'b101000000101101010111101111100000001000011000000010011,
        //tile 12
        54'b101000111101111100000101101010000001000011000000000000,
        //tile 13
        54'b101000111100111101000101101010000001000011000000000001,
        //tile 14
        54'b101000111101000101101010111100000001000011000000000010,
        //tile 15
        54'b101000000101101010111101111100000001000011000000000011,
        //tile 16
        54'b101000111101111100000101101010000001000011000000001100,
        //tile 17
        54'b101000111100111101000101101010000001000011000000001101,
        //tile 18
        54'b101000111101000101101010111100000001000011000000001110,
        //tile 19
        54'b101000000101101010111101111100000001000011000000001111,
        //tile 20
        54'b101000111101111100000101101010000001000011000000000000,
        //tile 21
        54'b101000111100111101000101101010000001000011000000000001,
        //tile 22
        54'b101000111101000101101010111100000001000011000000000010,
        //tile 23
        54'b101000000101101010111101111100000001000011000000000011,
        //tile 24
        54'b101000111101111100000101101010000001000011000000010000,
        //tile 25
        54'b101000111100111101000101101010000001000011000000010001,
        //tile 26
        54'b101000111101000101101010111100000001000011000000010010,
        //tile 27
        54'b101000000101101010111101111100000001000011000000010011,
        //tile 28
        54'b101000111101111100000101101010000001000011000000000000,
        //tile 29
        54'b101000111100111101000101101010000001000011000000000001,
        //tile 30
        54'b101000111101000101101010111100000001000011000000000010,
        //tile 31
        54'b101000000101101010111101111100000001000011000000000011,

        // <--- FILE: ASSETS\PLAYER\3-DEATH.PNG --->

        //tile 0
        54'b101000111101111100000101101010000001000011000000000000,
        //tile 1
        54'b101000111100111101000101101010000001000011000000000001,
        //tile 2
        54'b101000111101000101101010111100000001000011000000000010,
        //tile 3
        54'b101000000101101010111101111100000001000011000000000011,
        //tile 4
        54'b101000111101111100000101101010000001000011000000000000,
        //tile 5
        54'b101000111100111101000101101010000001000011000000000001,
        //tile 6
        54'b101000111101000101101010111100000001000011000000000010,
        //tile 7
        54'b101000000101101010111101111100000001000011000000000011,
        //tile 8
        54'b101000111101111100000101111110000001000011000000010100,
        //tile 9
        54'b101000111100111101000101111110000001000011000000010101,
        //tile 10
        54'b101000111101000101111110111100000001000011000000010110,
        //tile 11
        54'b101000000101111110111101111100000001000011000000010111,
        //tile 12
        54'b101000111101111100000101111110000001000011000000010100,
        //tile 13
        54'b101000111100111101000101111110000001000011000000011000,
        //tile 14
        54'b101000111101000101111110111100000001000011000000011001,
        //tile 15
        54'b101000000101111110111101111100000001000011000000011010,
        //tile 16
        54'b101000111101111100000101101010000001000011000000000000,
        //tile 17
        54'b101000111100111101000101101010000001000011000000000001,
        //tile 18
        54'b101000111101000101101010111100000001000011000000000010,
        //tile 19
        54'b101000000101101010111101111100000001000011000000000011,
        //tile 20
        54'b101000111101111100000101101010000001000011000000000000,
        //tile 21
        54'b101000111100111101000101101010000001000011000000000001,
        //tile 22
        54'b101000111101000101101010111100000001000011000000000010,
        //tile 23
        54'b101000000101101010111101111100000001000011000000000011,
        //tile 24
        54'b101000111101111100000101111110000001000011000000010100,
        //tile 25
        54'b101000111100111101000101111110000001000011000000011000,
        //tile 26
        54'b101000111101000101111110111100000001000011000000011001,
        //tile 27
        54'b101000000101111110111101111100000001000011000000011010,
        //tile 28
        54'b101000111101111100000101111110000001000011000000010100,
        //tile 29
        54'b101000111100111101000101111110000001000011000000011000,
        //tile 30
        54'b101000111101000101111110111100000001000011000000011001,
        //tile 31
        54'b101000000101111110111101111100000001000011000000011010,
        //tile 32
        54'b000000000000000000111101111100000001000011000000011011,
        //tile 33
        54'b000000000000000000111100111101000001000011000000011100,
        //tile 34
        54'b000000000000000000111101111100000001000011000000011101,
        //tile 35
        54'b000000000000000000111101111100000001000011000000011110,
        //tile 36
        54'b000000000000000000111101111100000001000011000000011111,
        //tile 37
        54'b000000000000000000111100111101000001000011000000100000,
        //tile 38
        54'b000000000000000000111100111101000001000011000000100001,
        //tile 39
        54'b000000000000000000111101111100000001000011000000100010,
        //tile 40
        54'b000000000000000000000000000001000011111101000000100011,
        //tile 41
        54'b000000000000000000000001000011111100111101000000100100,
        //tile 42
        54'b000000000000000000000000000001000011111101000000100101,
        //tile 43
        54'b000000000000000000000001000011111100111101000000100110,
        //tile 44
        54'b000000000000000000000001000011111100111101000000100111,
        //tile 45
        54'b000000000000000000000001000011111100111101000000101000,
        //tile 46
        54'b000000000000000000000001000011111100111101000000101001,
        //tile 47
        54'b000000000000000000000001000011111100111101000000101010,
        //tile 48
        54'b000000000000000000000001000011111100111101000000100111,
        //tile 49
        54'b000000000000000000000001000011111100111101000000101000,
        //tile 50
        54'b000000000000000000000001000011111100111101000000101001,
        //tile 51
        54'b000000000000000000000001000011111100111101000000101010,
        //tile 52
        54'b000000000000000000000001000011111100111101000000100111,
        //tile 53
        54'b000000000000000000000001000011111100111101000000101000,
        //tile 54
        54'b000000000000000000000001000011111100111101000000101001,
        //tile 55
        54'b000000000000000000000001000011111100111101000000101010,
        //tile 56
        54'b000000000000000000000001000011111100111101000000100111,
        //tile 57
        54'b000000000000000000000001000011111100111101000000101000,
        //tile 58
        54'b000000000000000000000001000011111100111101000000101001,
        //tile 59
        54'b000000000000000000000001000011111100111101000000101010,
        //tile 60
        54'b000000000000000000000001000011111100111101000000100111,
        //tile 61
        54'b000000000000000000000001000011111100111101000000101000,
        //tile 62
        54'b000000000000000000000001000011111100111101000000101001,
        //tile 63
        54'b000000000000000000000001000011111100111101000000101010
    
    };

    localparam bit [95:0] BITMAPS [1376] = '{


        // <--- FILE: ASSETS\PLAYER\1-IDLE.PNG --->

        //tile 0, VRAM 54'b101000111101111100000101101010000001000011000000000000
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000101101110011011011011011011011011011011011011011000000000,
        96'b000000000000000000000000000000000000000101101110011011011011011011011011011011011011011000000000,
        96'b000000000000000000000000000000101101101110110110101011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000101101101110110110110011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000101110110110110110110110101101101011011011011011011011000000000000,
        96'b000000000000000000000000000000101110110110110110110110110110101011011011011011011011000000000000,
        96'b000000000000000000000000000000110110110110110110110011011011011111111111111111111111000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011111111111111111111111000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        //tile 1, VRAM 54'b101000111100111101000101101010000001000011000000000001
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000101101101101110110110011011011011011011011011011011011011011000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011011000000000,
        96'b000000000000000000000101101101101101101101101101110011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101110101101101101101011011011011011011011011011011011000000000000,
        96'b000000000000000000101101101110110101101101101101101101110110110011011011011011011011000000000000,
        96'b000000000000000000101101101101101101101101101101101101101101110011011011011011011011000000000000,
        96'b000000000000000000101101101101101101101101101101101011011011011111111111111111111111000000000000,
        96'b000000000000000000101101101101101101101101101101011011011011011111111111111111111111000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        //tile 2, VRAM 54'b101000111101000101101010111100000001000011000000000010
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000011011011011000000100100100100100101101010100101010010100000000000,
        96'b000000000000000000000000011011110110110110011011100100100100100101101010100101010010100000000000,
        96'b000000000000000110110110110110110110110110110110100100100100100100100100100100100100100000000000,
        96'b000000000000000110110110110110110110110110110110100100100100100100100100100100100100100000000000,
        96'b000000000000110110110110110110110110110110110110011100100100100100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110100100100100100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110110011011011100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110110110110011100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110100100100100111111111111111111111000000000000,
        96'b000000000000110110110110110110110110110110110110100100100100100111111111111111111111000000000000,
        96'b000000000000110110110110110110110110011011110110100100100100100100100100100100100100000000000000,
        96'b000000000000011110110110110110011011110110110110100100100100100100100100100100100100000000000000,
        96'b000000000000000011011110110110110110110110110110100100100100100100100100100100100100000000000000,
        96'b000000000000000000000110110110110110110110110110100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100000000000100100100100100100000,
        96'b000000000000000000000000000000000000000000000000100100100100100100000000000100100100100100100000,
        //tile 3, VRAM 54'b101000000101101010111101111100000001000011000000000011
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000011011011011011011011011000001001001001001001001001001001001001001001001001,
        96'b000000000000000000011011100100100011011011011011101101101101101110110010101110010010101000000000,
        96'b000000000000000011100100100100100100100100100011101101101101101110110010101110010010101000000000,
        96'b000000000011011100100100100100100100100100100011101101101101101101101101101101101101101000000000,
        96'b000000100100100100100100100100100100100100100100101101101101101101101101101101101101101000000000,
        96'b000000100100100100100100100100100100100100100100011101101101101101101101101101101101000000000000,
        96'b000100100100100100100100100100100100100100100100100101101101101101101101101101101101000000000000,
        96'b000100100100100100011100100100100100100100100100100100011011011101101101101101101101000000000000,
        96'b000100100100100100011100100100100100100100100100100100100100011101101101101101101101000000000000,
        96'b000100100100100100011011100100100100100100100100100101101101101111111111111111111111000000000000,
        96'b000100100100100100100011100100100100100100100100101101101101101111111111111111111111000000000000,
        96'b000100100100100100100011011011100100100100100100101101101101101101101101101101101101000000000000,
        96'b000100100100100100100100100011011100100100100100101101101101101101101101101101101101000000000000,
        96'b000100100100100100100100100100100100100100100100101101101101101101101101101101101101000000000000,
        96'b000000100100100100100100100100100100100100100100101101101101101101101101101101101101000000000000,
        96'b000000000100100100100100100100100100100100100100101101101101101101101101101101101101000000000000,
        96'b000000000000000100100100100100100100100100000000101101101101101101101101101101101101000000000000,
        96'b000000000000000000000100100100100100000000000000101101101101101101101101101101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101000000000000000000101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101000000000000000000101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101000000000000000000101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101000000000000000000101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101101101101000000000101101101101101101000,
        96'b000000000000000000000000000000000000000000000000101101101101101101000000000101101101101101101000,
        //tile 4, VRAM 54'b101000111101111100000101101010000001000011000000000100
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000101101110011011011011011011011011011011011011011000000000,
        96'b000000000000000000000000000000000000000101101110101011011011011011011011011011011011011000000000,
        96'b000000000000000000000000000000101101101110110110110011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000101101101110110110110110101101101011011011011011011011000000000000,
        96'b000000000000000000000000000000101110110110110110110110110110101011011011011011011011000000000000,
        96'b000000000000000000000000000000101110110110110110110110110110101011011011011011011011000000000000,
        96'b000000000000000000000000000000110110110110110110110011011011011111111111111111111111000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011111111111111111111111000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        //tile 5, VRAM 54'b101000111100111101000101101010000001000011000000000101
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000101101101101110110110011011011011011011011011011011011011011000000000,
        96'b000000000000000000000101101101101101101101101101110011011011011011011011011011011011011000000000,
        96'b000000000000000000000101101101101101101101101101101011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101110101101101101101101110110110011011011011011011011000000000000,
        96'b000000000000000000101101101110110101101101101101101101101101110011011011011011011011000000000000,
        96'b000000000000000000101101101101101101101101101101101101101101110011011011011011011011000000000000,
        96'b000000000000000000101101101101101101101101101101101011011011011111111111111111111111000000000000,
        96'b000000000000000000101101101101101101101101101101011011011011011111111111111111111111000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        //tile 6, VRAM 54'b101000111101111100000101101010000001000011000000000110
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000101101101101000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000101101110110110110101101011011011011011100100010011100010010011000000000,
        96'b000000000000000110110110110110110110110110110110011011011011011011011011011011011011011000000000,
        96'b000000000000000110110110110110110110110110110110101011011011011011011011011011011011011000000000,
        96'b000000000000110110110110110110110110110110110110110011011011011011011011011011011011000000000000,
        96'b000000000000110110110110110110110110110110110110110110101101101011011011011011011011000000000000,
        96'b000000000000110110110110110110110110110110110110110110110110101011011011011011011011000000000000,
        96'b000000000000110110110110110110110110110110110110110110110110101011011011011011011011000000000000,
        96'b000000000000110110110110110110110110110110110110110011011011011111111111111111111111000000000000,
        96'b000000000000110110110110110110110110110110110110011011011011011111111111111111111111000000000000,
        96'b000000000000110110110110110110110110101101110110011011011011011011011011011011011011000000000000,
        96'b000000000000101110110110110110101101110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000101101110110110110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000110110110110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        //tile 7, VRAM 54'b101000111101000101101010111100000001000011000000000111
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000011011011011011011011011000100100100100100101101010100101010010100000000000,
        96'b000000000000000000011011110110110011011011011011100100100100100101101010100101010010100000000000,
        96'b000000000000000011110110110110110110110110110011100100100100100101101010100101010010100000000000,
        96'b000000000011011110110110110110110110110110110011100100100100100100100100100100100100100000000000,
        96'b000000110110110110110110110110110110110110110110011100100100100100100100100100100100100000000000,
        96'b000000110110110110110110110110110110110110110110110100100100100100100100100100100100000000000000,
        96'b000110110110110110110110110110110110110110110110110110011011011100100100100100100100000000000000,
        96'b000110110110110110011110110110110110110110110110110110110110011100100100100100100100000000000000,
        96'b000110110110110110011110110110110110110110110110110110110110011100100100100100100100000000000000,
        96'b000110110110110110011011110110110110110110110110110100100100100111111111111111111111000000000000,
        96'b000110110110110110110011110110110110110110110110100100100100100111111111111111111111000000000000,
        96'b000110110110110110110011011011110110110110110110100100100100100100100100100100100100000000000000,
        96'b000110110110110110110110110011011110110110110110100100100100100100100100100100100100000000000000,
        96'b000110110110110110110110110110110110110110110110100100100100100100100100100100100100000000000000,
        96'b000000110110110110110110110110110110110110110110100100100100100100100100100100100100000000000000,
        96'b000000000110110110110110110110110110110110110110100100100100100100100100100100100100000000000000,
        96'b000000000000000110110110110110110110110110000000100100100100100100100100100100100100000000000000,
        96'b000000000000000000000110110110110110000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100000000000100100100100100100000,
        96'b000000000000000000000000000000000000000000000000100100100100100100000000000100100100100100100000,
        //tile 8, VRAM 54'b101000111101111100000101101010000001000011000000001000
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000101101110011011011011011011011011011011011011011000000000,
        96'b000000000000000000000000000000000000000101101110101011011011011011011011011011011011011000000000,
        96'b000000000000000000000000000000101101101110110110110011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000101101101110110110110110101101101011011011011011011011000000000000,
        96'b000000000000000000000000000000101110110110110110110110110110101011011011011011011011000000000000,
        96'b000000000000000000000000000000101110110110110110110110110110101011011011011011011011000000000000,
        96'b000000000000000000000000000000110110110110110110110011011011011111111111111111111111000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011111111111111111111111000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        //tile 9, VRAM 54'b101000111100111101000101101010000001000011000000001001
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000101101101101110110110011011011011011011011011011011011011011000000000,
        96'b000000000000000000000101101101101101101101101101110011011011011011011011011011011011011000000000,
        96'b000000000000000000000101101101101101101101101101101011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101110101101101101101101110110110011011011011011011011000000000000,
        96'b000000000000000000101101101110110101101101101101101101101101110011011011011011011011000000000000,
        96'b000000000000000000101101101101101101101101101101101101101101110011011011011011011011000000000000,
        96'b000000000000000000101101101101101101101101101101101011011011011111111111111111111111000000000000,
        96'b000000000000000000101101101101101101101101101101011011011011011111111111111111111111000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        //tile 10, VRAM 54'b101000111101111100000101101010000001000011000000001010
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000101101101101000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000101101110110110110101101011011011011011100100010011100010010011000000000,
        96'b000000000000000110110110110110110110110110110110011011011011011011011011011011011011011000000000,
        96'b000000000000000110110110110110110110110110110110101011011011011011011011011011011011011000000000,
        96'b000000000000110110110110110110110110110110110110110011011011011011011011011011011011000000000000,
        96'b000000000000110110110110110110110110110110110110110110101101101011011011011011011011000000000000,
        96'b000000000000110110110110110110110110110110110110110110110110101011011011011011011011000000000000,
        96'b000000000000110110110110110110110110110110110110110110110110101011011011011011011011000000000000,
        96'b000000000000110110110110110110110110110110110110110011011011011111111111111111111111000000000000,
        96'b000000000000110110110110110110110110110110110110011011011011011111111111111111111111000000000000,
        96'b000000000000110110110110110110110110101101110110011011011011011011011011011011011011000000000000,
        96'b000000000000101110110110110110101101110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000101101110110110110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000110110110110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        //tile 11, VRAM 54'b101000111101000101101010111100000001000011000000001011
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000011011011011011011011011000100100100100100101101010100101010010100000000000,
        96'b000000000000000000011011110110110011011011011011100100100100100101101010100101010010100000000000,
        96'b000000000000000011110110110110110110110110110011100100100100100101101010100101010010100000000000,
        96'b000000000011011110110110110110110110110110110011100100100100100100100100100100100100100000000000,
        96'b000000110110110110110110110110110110110110110110011100100100100100100100100100100100100000000000,
        96'b000000110110110110110110110110110110110110110110110100100100100100100100100100100100000000000000,
        96'b000110110110110110110110110110110110110110110110110110011011011100100100100100100100000000000000,
        96'b000110110110110110011110110110110110110110110110110110110110011100100100100100100100000000000000,
        96'b000110110110110110011110110110110110110110110110110110110110011100100100100100100100000000000000,
        96'b000110110110110110011011110110110110110110110110110100100100100111111111111111111111000000000000,
        96'b000110110110110110110011110110110110110110110110100100100100100111111111111111111111000000000000,
        96'b000110110110110110110011011011110110110110110110100100100100100100100100100100100100000000000000,
        96'b000110110110110110110110110011011110110110110110100100100100100100100100100100100100000000000000,
        96'b000110110110110110110110110110110110110110110110100100100100100100100100100100100100000000000000,
        96'b000000110110110110110110110110110110110110110110100100100100100100100100100100100100000000000000,
        96'b000000000110110110110110110110110110110110110110100100100100100100100100100100100100000000000000,
        96'b000000000000000110110110110110110110110110000000100100100100100100100100100100100100000000000000,
        96'b000000000000000000000110110110110110000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100000000000100100100100100100000,
        96'b000000000000000000000000000000000000000000000000100100100100100100000000000100100100100100100000,

        // <--- FILE: ASSETS\PLAYER\2-WALK.PNG --->

        //tile 12, VRAM 54'b101000111101111100000101101010000001000011000000001100
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000101101110011011011011011011011011011011011011011000000000,
        96'b000000000000000000000000000000000000000101101110011011011011011011011011011011011011011000000000,
        96'b000000000000000000000000000000101101101110110110101011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000101101101110110110110011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000101110110110110110110110101101101011011011011011011011000000000000,
        96'b000000000000000000000000000000101110110110110110110110110110101011011011011011011011000000000000,
        96'b000000000000000000000000000000110110110110110110110011011011011111111111111111111111000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011111111111111111111111000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000,
        //tile 13, VRAM 54'b101000111100111101000101101010000001000011000000001101
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000101101101101110110110011011011011011011011011011011011011011000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011011000000000,
        96'b000000000000000000000101101101101101101101101101110011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101110101101101101101011011011011011011011011011011011000000000000,
        96'b000000000000000000101101101110110101101101101101101101110110110011011011011011011011000000000000,
        96'b000000000000000000101101101101101101101101101101101101101101110011011011011011011011000000000000,
        96'b000000000000000000101101101101101101101101101101101011011011011111111111111111111111000000000000,
        96'b000000000000000000101101101101101101101101101101011011011011011111111111111111111111000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000000000000000000000000,
        //tile 14, VRAM 54'b101000111101000101101010111100000001000011000000001110
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000011011011011000000100100100100100101101010100101010010100000000000,
        96'b000000000000000000000000011011110110110110011011100100100100100101101010100101010010100000000000,
        96'b000000000000000110110110110110110110110110110110100100100100100100100100100100100100100000000000,
        96'b000000000000000110110110110110110110110110110110100100100100100100100100100100100100100000000000,
        96'b000000000000110110110110110110110110110110110110011100100100100100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110100100100100100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110110011011011100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110110110110011100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110100100100100111111111111111111111000000000000,
        96'b000000000000110110110110110110110110110110110110100100100100100111111111111111111111000000000000,
        96'b000000000000110110110110110110110110011011110110100100100100100100100100100100100100000000000000,
        96'b000000000000011110110110110110011011110110110110100100100100100100100100100100100100000000000000,
        96'b000000000000000011011110110110110110110110110110100100100100100100100100100100100100000000000000,
        96'b000000000000000000000110110110110110110110110110100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100100100100000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100100100100000,
        96'b000000000000000000000000000000000000000000000000100100100100100100000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100000000000000000000000000000000,
        //tile 15, VRAM 54'b101000000101101010111101111100000001000011000000001111
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000011011011011011011011011000001001001001001001001001001001001001001001001001,
        96'b000000000000000000011011100100100011011011011011101101101101101110110010101110010010101000000000,
        96'b000000000000000011100100100100100100100100100011101101101101101110110010101110010010101000000000,
        96'b000000000011011100100100100100100100100100100011101101101101101101101101101101101101101000000000,
        96'b000000100100100100100100100100100100100100100100101101101101101101101101101101101101101000000000,
        96'b000000100100100100100100100100100100100100100100011101101101101101101101101101101101000000000000,
        96'b000100100100100100100100100100100100100100100100100101101101101101101101101101101101000000000000,
        96'b000100100100100100011100100100100100100100100100100100011011011101101101101101101101000000000000,
        96'b000100100100100100011100100100100100100100100100100100100100011101101101101101101101000000000000,
        96'b000100100100100100011011100100100100100100100100100101101101101111111111111111111111000000000000,
        96'b000100100100100100100011100100100100100100100100101101101101101111111111111111111111000000000000,
        96'b000100100100100100100011011011100100100100100100101101101101101101101101101101101101000000000000,
        96'b000100100100100100100100100011011100100100100100101101101101101101101101101101101101000000000000,
        96'b000100100100100100100100100100100100100100100100101101101101101101101101101101101101000000000000,
        96'b000000100100100100100100100100100100100100100100101101101101101101101101101101101101000000000000,
        96'b000000000100100100100100100100100100100100100100101101101101101101101101101101101101000000000000,
        96'b000000000000000100100100100100100100100100000000101101101101101101101101101101101101000000000000,
        96'b000000000000000000000100100100100100000000000000101101101101101101101101101101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101000000000000000000101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101000000000000000000101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101000000000000000000101101101101101101000,
        96'b000000000000000000000000000000000000000000000000101101101000000000000000000101101101101101101000,
        96'b000000000000000000000000000000000000000000000000101101101101101101000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000101101101101101101000000000000000000000000000000,
        //tile 16, VRAM 54'b101000111101111100000101101010000001000011000000010000
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000000,
        96'b000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000000,
        96'b000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000,
        96'b000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000,
        96'b000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000,
        96'b000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000000,
        96'b000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000000,
        96'b000000000000000000000000000000000000101101110011011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000101101110011011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000101101101110110110101011011011011011011011011011011011000000000000000,
        96'b000000000000000000000000000101101101110110110110011011011011011011011011011011011000000000000000,
        96'b000000000000000000000000000101110110110110110110110101101101011011011011011011011000000000000000,
        96'b000000000000000000000000000101110110110110110110110110110101011011011011011011011000000000000000,
        96'b000000000000000000000000000110110110110110110110011011011011111111111111111111111000000000000000,
        96'b000000000000000000000000000110110110110110110011011011011011111111111111111111111000000000000000,
        96'b000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000000,
        96'b000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000000,
        96'b000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000000,
        96'b000000000000000000000000000000110110110110110011011011011011011011011011011011011000000000000000,
        96'b000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        96'b000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        96'b000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        96'b000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000000,
        96'b000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000000,
        96'b000000000000000000000000000000000000000000000011011011011011011000000000011011011000000000000000,
        96'b000000000000000000000000000000000000000000000011011011011011011000000000011011011000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011000000,
        //tile 17, VRAM 54'b101000111100111101000101101010000001000011000000010001
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000000,
        96'b000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000000,
        96'b000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000,
        96'b000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000,
        96'b000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000,
        96'b000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000000,
        96'b000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000000,
        96'b000000000000000000000000101101101101110110110011011011011011011011011011011011011011000000000000,
        96'b000000000000000000101101101101101101101101101011011011011011011011011011011011011011000000000000,
        96'b000000000000000000101101101101101101101101101110011011011011011011011011011011011000000000000000,
        96'b000000000000000000101101101101110101101101101101011011011011011011011011011011011000000000000000,
        96'b000000000000000101101101110110101101101101101101101110110110011011011011011011011000000000000000,
        96'b000000000000000101101101101101101101101101101101101101101110011011011011011011011000000000000000,
        96'b000000000000000101101101101101101101101101101101011011011011111111111111111111111000000000000000,
        96'b000000000000000101101101101101101101101101101011011011011011111111111111111111111000000000000000,
        96'b000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000000,
        96'b000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000000,
        96'b000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000000,
        96'b000000000000000000000000101101101101101101101011011011011011011011011011011011011000000000000000,
        96'b000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        96'b000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        96'b000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000000,
        96'b000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000000,
        96'b000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000000,
        96'b000000000000000000000000000000000000000000000011011011011011011000000000011011011000000000000000,
        96'b000000000000000000000000000000000000000000000011011011011011011000000000011011011000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011000000,
        //tile 18, VRAM 54'b101000111101000101101010111100000001000011000000010010
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000000,
        96'b000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000000,
        96'b000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000,
        96'b000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000,
        96'b000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001000,
        96'b000000000000000000000000000011011011011000000100100100100100101101010100101010010100000000000000,
        96'b000000000000000000000011011110110110110011011100100100100100101101010100101010010100000000000000,
        96'b000000000000110110110110110110110110110110110100100100100100100100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110100100100100100100100100100100100100100000000000000,
        96'b000000000110110110110110110110110110110110110011100100100100100100100100100100100000000000000000,
        96'b000000000110110110110110110110110110110110110110100100100100100100100100100100100000000000000000,
        96'b000000000110110110110110110110110110110110110110110011011011100100100100100100100000000000000000,
        96'b000000000110110110110110110110110110110110110110110110110011100100100100100100100000000000000000,
        96'b000000000110110110110110110110110110110110110110100100100100111111111111111111111000000000000000,
        96'b000000000110110110110110110110110110110110110100100100100100111111111111111111111000000000000000,
        96'b000000000110110110110110110110110011011110110100100100100100100100100100100100100000000000000000,
        96'b000000000011110110110110110011011110110110110100100100100100100100100100100100100000000000000000,
        96'b000000000000011011110110110110110110110110110100100100100100100100100100100100100000000000000000,
        96'b000000000000000000110110110110110110110110110100100100100100100100100100100100100000000000000000,
        96'b000000000000000000000000000000000000000000000100100100100100100100100100100100100000000000000000,
        96'b000000000000000000000000000000000000000000000100100100100100100100100100100100100000000000000000,
        96'b000000000000000000000000000000000000000000000100100100100100100100100100100100100000000000000000,
        96'b000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000000,
        96'b000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000000,
        96'b000000000000000000000000000000000000000000000100100100100100100000000000100100100000000000000000,
        96'b000000000000000000000000000000000000000000000100100100100100100000000000100100100000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000100100100100100100000000,
        //tile 19, VRAM 54'b101000000101101010111101111100000001000011000000010011
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000000,
        96'b000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000000,
        96'b000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001001,
        96'b000000000000000000011011011011011011011011000001001001001001001001001001001001001001001001001001,
        96'b000000000000000011011100100100011011011011011101101101101101110110010101110010010101000000000000,
        96'b000000000000011100100100100100100100100100011101101101101101110110010101110010010101000000000000,
        96'b000000011011100100100100100100100100100100011101101101101101101101101101101101101101000000000000,
        96'b000100100100100100100100100100100100100100100101101101101101101101101101101101101101000000000000,
        96'b000100100100100100100100100100100100100100100011101101101101101101101101101101101000000000000000,
        96'b100100100100100100100100100100100100100100100100101101101101101101101101101101101000000000000000,
        96'b100100100100100011100100100100100100100100100100100011011011101101101101101101101000000000000000,
        96'b100100100100100011100100100100100100100100100100100100100011101101101101101101101000000000000000,
        96'b100100100100100011011100100100100100100100100100101101101101111111111111111111111000000000000000,
        96'b100100100100100100011100100100100100100100100101101101101101111111111111111111111000000000000000,
        96'b100100100100100100011011011100100100100100100101101101101101101101101101101101101000000000000000,
        96'b100100100100100100100100011011100100100100100101101101101101101101101101101101101000000000000000,
        96'b100100100100100100100100100100100100100100100101101101101101101101101101101101101000000000000000,
        96'b000100100100100100100100100100100100100100100101101101101101101101101101101101101000000000000000,
        96'b000000100100100100100100100100100100100100100101101101101101101101101101101101101000000000000000,
        96'b000000000000100100100100100100100100100000000101101101101101101101101101101101101000000000000000,
        96'b000000000000000000100100100100100000000000000101101101101101101101101101101101101000000000000000,
        96'b000000000000000000000000000000000000000000000101101101000000000000000000101101101000000000000000,
        96'b000000000000000000000000000000000000000000000101101101000000000000000000101101101000000000000000,
        96'b000000000000000000000000000000000000000000000101101101101101101000000000101101101000000000000000,
        96'b000000000000000000000000000000000000000000000101101101101101101000000000101101101000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000101101101101101101000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000101101101101101101000000,

        // <--- FILE: ASSETS\PLAYER\3-DEATH.PNG --->

        //tile 20, VRAM 54'b101000111101111100000101111110000001000011000000010100
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000101101110011011011011011011011011011011011011011000000000,
        96'b000000000000000000000000000000000000000101101110011011011011011011011011011011011011011000000000,
        96'b000000000000000000000000000000101101101110110110101011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000101101101110110110110011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000101110110110110110110110101101101011011011011011011011000000000000,
        96'b000000000000000000000000000000101110110110110110110110110110101011011011011011011011000000000000,
        96'b000000000000000000000000000000110110110110110110110011011011011111111111111111111111000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011111111111111111111111000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000110110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000110110110110110011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        //tile 21, VRAM 54'b101000111100111101000101111110000001000011000000010101
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000101101101101110110110011011011011011011011011011011011011011000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011011000000000,
        96'b000000000000000000000101101101101101101101101101110011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101110101101101101101011011011011011011011011011011011000000000000,
        96'b000000000000000000101101101110110101101101101101101101110110110011011011011011011011000000000000,
        96'b000000000000000000101101101101101101101101101101101101101101110011011011011011011011000000000000,
        96'b000000000000000000101101101101101101101101101101101011011011011111111111111111111111000000000000,
        96'b000000000000000000101101101101101101101101101101011011011011011111111111111111111111000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        //tile 22, VRAM 54'b101000111101000101111110111100000001000011000000010110
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000011011011011000000100100100100100101101010100101010010100000000000,
        96'b000000000000000000000000011011110110110110011011100100100100100101101010100101010010100000000000,
        96'b000000000000000110110110110110110110110110110110100100100100100100100100100100100100100000000000,
        96'b000000000000000110110110110110110110110110110110100100100100100100100100100100100100100000000000,
        96'b000000000000110110110110110110110110110110110110011100100100100100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110100100100100100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110110011011011100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110110110110011100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110100100100100111111111111111111111000000000000,
        96'b000000000000110110110110110110110110110110110110100100100100100111111111111111111111000000000000,
        96'b000000000000110110110110110110110110011011110110100100100100100100100100100100100100000000000000,
        96'b000000000000011110110110110110011011110110110110100100100100100100100100100100100100000000000000,
        96'b000000000000000011011110110110110110110110110110100100100100100100100100100100100100000000000000,
        96'b000000000000000000000110110110110110110110110110100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100000000000100100100100100100000,
        96'b000000000000000000000000000000000000000000000000100100100100100100000000000100100100100100100000,
        //tile 23, VRAM 54'b101000000101111110111101111100000001000011000000010111
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000011011011011011011011011000001001001001001001001001001001001001001001001001,
        96'b000000000000000000011011100100100011011011011011101101101101101110110010101110010010101000000000,
        96'b000000000000000011100100100100100100100100100011101101101101101110110010101110010010101000000000,
        96'b000000000011011100100100100100100100100100100011101101101101101101101101101101101101101000000000,
        96'b000000100100100100100100100100100100100100100100101101101101101101101101101101101101101000000000,
        96'b000000100100100100100100100100100100100100100100011101101101101101101101101101101101000000000000,
        96'b000100100100100100100100100100100100100100100100100101101101101101101101101101101101000000000000,
        96'b000100100100100100011100100100100100100100100100100100011011011101101101101101101101000000000000,
        96'b000100100100100100011100100100100100100100100100100100100100011101101101101101101101000000000000,
        96'b000100100100100100011011100100100100100100100100100101101101101111111111111111111111000000000000,
        96'b000100100100100100100011100100100100100100100100101101101101101111111111111111111111000000000000,
        96'b000100100100100100100011011011100100100100100100101101101101101101101101101101101101000000000000,
        96'b000100100100100100100100100011011100100100100100101101101101101101101101101101101101000000000000,
        96'b000100100100100100100100100100100100100100100100101101101101101101101101101101101101000000000000,
        96'b000000100100100100100100100100100100100100100100101101101101101101101101101101101101000000000000,
        96'b000000000100100100100100100100100100100100100100101101101101101101101101101101101101000000000000,
        96'b000000000000000100100100100100100100100100000000101101101101101101101101101101101101000000000000,
        96'b000000000000000000000100100100100100000000000000101101101101101101101101101101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101000000000000000000101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101000000000000000000101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101000000000000000000101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101000000000000000000101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101101101101000000000101101101101101101000,
        96'b000000000000000000000000000000000000000000000000101101101101101101000000000101101101101101101000,
        //tile 24, VRAM 54'b101000111100111101000101111110000001000011000000011000
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011100100010011100010010011000000000,
        96'b000000000000000000000000000101101101101110110110011011011011011011011011011011011011011000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011011000000000,
        96'b000000000000000000000101101101101101101101101101110011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101110101101101101101011011011011011011011011011011011000000000000,
        96'b000000000000000000101101101110110101101101101101101101110110110011011011011011011011000000000000,
        96'b000000000000000000101101101101101101101101101101101101101101110011011011011011011011000000000000,
        96'b000000000000000000101101101101101101101101101101101011011011011111111111111111111111000000000000,
        96'b000000000000000000101101101101101101101101101101011011011011011111111111111111111111000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000101101101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000101101101101101101101011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011011011011011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011000000000000000000011011011000000000000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000011011011011011011000000000011011011011011011000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        //tile 25, VRAM 54'b101000111101000101111110111100000001000011000000011001
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000011011011011000000100100100100100101101010100101010010100000000000,
        96'b000000000000000000000000011011110110110110011011100100100100100101101010100101010010100000000000,
        96'b000000000000000110110110110110110110110110110110100100100100100100100100100100100100100000000000,
        96'b000000000000000110110110110110110110110110110110100100100100100100100100100100100100100000000000,
        96'b000000000000110110110110110110110110110110110110011100100100100100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110100100100100100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110110011011011100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110110110110011100100100100100100100000000000000,
        96'b000000000000110110110110110110110110110110110110110100100100100111111111111111111111000000000000,
        96'b000000000000110110110110110110110110110110110110100100100100100111111111111111111111000000000000,
        96'b000000000000110110110110110110110110011011110110100100100100100100100100100100100100000000000000,
        96'b000000000000011110110110110110011011110110110110100100100100100100100100100100100100000000000000,
        96'b000000000000000011011110110110110110110110110110100100100100100100100100100100100100000000000000,
        96'b000000000000000000000110110110110110110110110110100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100100100100100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100000000000000000000100100100000000000000,
        96'b000000000000000000000000000000000000000000000000100100100100100100000000000100100100100100100000,
        96'b000000000000000000000000000000000000000000000000100100100100100100000000000100100100100100100000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        //tile 26, VRAM 54'b101000000101111110111101111100000001000011000000011010
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000011011011011011011011011000001001001001001001001001001001001001001001001001,
        96'b000000000000000000011011100100100011011011011011101101101101101110110010101110010010101000000000,
        96'b000000000000000011100100100100100100100100100011101101101101101110110010101110010010101000000000,
        96'b000000000011011100100100100100100100100100100011101101101101101101101101101101101101101000000000,
        96'b000000100100100100100100100100100100100100100100101101101101101101101101101101101101101000000000,
        96'b000000100100100100100100100100100100100100100100011101101101101101101101101101101101000000000000,
        96'b000100100100100100100100100100100100100100100100100101101101101101101101101101101101000000000000,
        96'b000100100100100100011100100100100100100100100100100100011011011101101101101101101101000000000000,
        96'b000100100100100100011100100100100100100100100100100100100100011101101101101101101101000000000000,
        96'b000100100100100100011011100100100100100100100100100101101101101111111111111111111111000000000000,
        96'b000100100100100100100011100100100100100100100100101101101101101111111111111111111111000000000000,
        96'b000100100100100100100011011011100100100100100100101101101101101101101101101101101101000000000000,
        96'b000100100100100100100100100011011100100100100100101101101101101101101101101101101101000000000000,
        96'b000100100100100100100100100100100100100100100100101101101101101101101101101101101101000000000000,
        96'b000000100100100100100100100100100100100100100100101101101101101101101101101101101101000000000000,
        96'b000000000100100100100100100100100100100100100100101101101101101101101101101101101101000000000000,
        96'b000000000000000100100100100100100100100100000000101101101101101101101101101101101101000000000000,
        96'b000000000000000000000100100100100100000000000000101101101101101101101101101101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101000000000000000000101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101000000000000000000101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101000000000000000000101101101000000000000,
        96'b000000000000000000000000000000000000000000000000101101101101101101000000000101101101101101101000,
        96'b000000000000000000000000000000000000000000000000101101101101101101000000000101101101101101101000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        //tile 27, VRAM 54'b000000000000000000111101111100000001000011000000011011
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000011011100000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000011011011011011100000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000011011011100100100100000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000011011011100100100100000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000011100100100100100100100000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000011100100100100100100100000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000100100100100100100100100000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000100100100100100100100100000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000100100100100100100100100000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000100100100100100100000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000100100100100100100000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000100100100100100000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        //tile 28, VRAM 54'b000000000000000000111100111101000001000011000000011100
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000000000000000000000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000000011011011011100100100000000000000000000000000000000000000000000000000,
        96'b000000000000000000000011011011011011011011011011000000000000000000000000000000000000000000000000,
        96'b000000000000000000000011011011011011011011011011100000000000000000000000000000000000000000000000,
        96'b000000000000000000011011011011011100011011011011011000000000000000000000000000000000000000000000,
        96'b000000000000000000011011011100100011011011011011011011100000000000000000000000000000000000000000,
        96'b000000000000000000011011011011011011011011011011011011011011000000000000000000000000000000000000,
        96'b000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000,
        96'b000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000,
        96'b000000000000000000000011011011011011011011011011011011000000000000000000000000000000000000000000,
        96'b000000000000000000000011011011011011011011011011011000000000000000000000000000000000000000000000,
        96'b000000000000000000000011011011011011011011011011000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000011011011011011011011000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        //tile 29, VRAM 54'b000000000000000000111101111100000001000011000000011101
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000000000000011011011011000000001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000011011011011011011011011001001001001001001001001001001001001001001001001,
        96'b000000000000000000000000011011100100100100011011001001001001001001001001001001001001001001001001,
        96'b000000000000000100100100100100100100100100100100000000000000000000000000000000000000000000000000,
        96'b000000000000100100100100100100100100100100100100000000000000000000000000000000000000000000000000,
        96'b000000000000100100100100100100100100100100100100011000000000000000000000000000000000000000000000,
        96'b000000000000100100100100100100100100100100100100100000000000000000000000000000000000000000000000,
        96'b000000000000100100100100100100100100100100100100100100011000000000000000000000000000000000000000,
        96'b000000000000100100100100100100100100100100100100100100100000000000000000000000000000000000000000,
        96'b000000000000100100100100100100100100100100100100100100000000000000000000000000000000000000000000,
        96'b000000000000100100100100100100100100100100100100100100000000000000000000000000000000000000000000,
        96'b000000000000100100100100100100100100011011100100100100000000000000000000000000000000000000000000,
        96'b000000000000011100100100100100011011100100100100100000000000000000000000000000000000000000000000,
        96'b000000000000000011011100100100100100100100100100000000000000000000000000000000000000000000000000,
        96'b000000000000000000000100100100100100100100100100000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        //tile 30, VRAM 54'b000000000000000000111101111100000001000011000000011110
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000001010010010010010010010010010010010010000000000,
        96'b000000000000000000000011011011011011011011011000001010010010010010010010010010010010010000000000,
        96'b000000000000000000011011011011011011011011011011001001001001001001001001001001001001001001001001,
        96'b000000000000000011011011100100100011011011011011001001001001001001001001001001001001001001001001,
        96'b000000000000000011100100100100100100100100100011001001001001001001001001001001001001001001001001,
        96'b000000000011011100100100100100100100100100100011000000000000000000000000000000000000000000000000,
        96'b000000100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000,
        96'b000100100100100100100100100100100100100100100100011000000000000000000000000000000000000000000000,
        96'b000100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000,
        96'b000100100100100100011100100100100100100100100100100100011000000000000000000000000000000000000000,
        96'b000100100100100100011100100100100100100100100100100100100100000000000000000000000000000000000000,
        96'b000100100100100100011011100100100100100100100100100100000000000000000000000000000000000000000000,
        96'b000100100100100100100011100100100100100100100100100100000000000000000000000000000000000000000000,
        96'b000100100100100100100011011011100100100100100100100100000000000000000000000000000000000000000000,
        96'b000100100100100100100100100011011100100100100100100000000000000000000000000000000000000000000000,
        96'b000100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000,
        96'b000000100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000,
        96'b000000000100100100100100100100100100100100100100000000000000000000000000000000000000000000000000,
        96'b000000000000000100100100100100100100100100000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000100100100100100000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        //tile 31, VRAM 54'b000000000000000000111101111100000001000011000000011111
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000001010010010010010010010010010010010010000000000000000000000000000000000000,
        96'b000000000000000000000001010010010010010010010010010010010010000000000000000000000000000000000000,
        96'b000000000000000000000001001001001001001001001001001001001001001001001000000000000000000000000000,
        96'b000000000000000000000001001001001001001001001001001001001001001001001000000000000000000000000000,
        96'b000000000000000000000001001001001001001001001001001001001001001001001000000000000000000000000000,
        96'b000000000000000000000000000000011011011100100100100000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000011100100100100100100100000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000011100100100100100100100000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000100100100100100100100100000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000100100100100100100100100000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000100100100100100100100100000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000100100100100100100000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000100100100100100100000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        //tile 32, VRAM 54'b000000000000000000111100111101000001000011000000100000
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000001010010010010010010010010010010010010000000000000000000000000000000000,
        96'b000000000000000000000000001010010010010010010010010010010010010000000000000000000000000000000000,
        96'b000000000000000000000000001001001001001001001001001001001001001001001001000000000000000000000000,
        96'b000000000000000000000000001001001001001001001001001001001001001001001001000000000000000000000000,
        96'b000000000000000000000011001001001001001001001001001001001001001001001001000000000000000000000000,
        96'b000000000000000000011011011011011100011011011011011000000000000000000000000000000000000000000000,
        96'b000000000000000000011011011100100011011011011011011011100000000000000000000000000000000000000000,
        96'b000000000000000000011011011011011011011011011011011011011000000000000000000000000000000000000000,
        96'b000000000000000000011011011011011011011011011011011011011000000000000000000000000000000000000000,
        96'b000000000000000000011011011011011011011011011011011011000000000000000000000000000000000000000000,
        96'b000000000000000000000011011011011011011011011011011000000000000000000000000000000000000000000000,
        96'b000000000000000000000011011011011011011011011011000000000000000000000000000000000000000000000000,
        96'b000000000000000000000011011011011011011011011011000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        //tile 33, VRAM 54'b000000000000000000111100111101000001000011000000100001
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000001010010010010010010010010010010010010000000000000000000000000000000000000,
        96'b000000000000000000000001010010010010010010010010010010010010000000000000000000000000000000000000,
        96'b000000000000000000000001001001001001001001001001001001001001001001001000000000000000000000000000,
        96'b000000000000000011011001001001001001001001001001001001001001001001001000000000000000000000000000,
        96'b000000000000011011011001001001001001001001001001001001001001001001001000000000000000000000000000,
        96'b000000000000011011011011011011011011011011011011011000000000000000000000000000000000000000000000,
        96'b000000000000011011011011011011011011011011011011011011100000000000000000000000000000000000000000,
        96'b000000000000011011011011011011011011011011011011011011011000000000000000000000000000000000000000,
        96'b000000000000011011011011011011011011011011011011011011011000000000000000000000000000000000000000,
        96'b000000000000011011011011011011011011011011011011011011000000000000000000000000000000000000000000,
        96'b000000000000011011011011011011011011100100011011011011000000000000000000000000000000000000000000,
        96'b000000000000100011011011011011100100011011011011011000000000000000000000000000000000000000000000,
        96'b000000000000000100100011011011011011011011011011000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        //tile 34, VRAM 54'b000000000000000000111101111100000001000011000000100010
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000001010010010010010010010010010010010010000000000000000000000000000000000,
        96'b000000000000000000000011001010010010010010010010010010010010010000000000000000000000000000000000,
        96'b000000000000000011100100001001001001001001001001001001001001001001001001000000000000000000000000,
        96'b000000000011011100100100001001001001001001001001001001001001001001001001000000000000000000000000,
        96'b000000100100100100100100001001001001001001001001001001001001001001001001000000000000000000000000,
        96'b000100100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000,
        96'b000100100100100100011100100100100100100100100100100100100000000000000000000000000000000000000000,
        96'b000100100100100100011100100100100100100100100100100100100000000000000000000000000000000000000000,
        96'b000100100100100100011011100100100100100100100100100100100000000000000000000000000000000000000000,
        96'b000100100100100100100011100100100100100100100100100100100000000000000000000000000000000000000000,
        96'b000100100100100100100011011011100100100100100100100100100000000000000000000000000000000000000000,
        96'b000100100100100100100100100011011100100100100100100100000000000000000000000000000000000000000000,
        96'b000100100100100100100100100100100100100100100100000000000000000000000000000000000000000000000000,
        96'b000000000000000100100100100100100100100100000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000100100100100100000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        //tile 35, VRAM 54'b000000000000000000000000000001000011111101000000100011
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000010011011011011011011011011011011011011000000000000000000000000000000,
        96'b000000000000000000000000000010011011011011011011011011011011011011000000000000000000000000000000,
        96'b000000000000000000000000000010010010010010010010010010010010010010010010010000000000000000000000,
        96'b000000000000000000000000000010010010010010010010010010010010010010010010010000000000000000000000,
        96'b000000000000000000000000000010010010010010010010010010010010010010010010010000000000000000000000,
        96'b000000000000000000000000000000001001001001001001001001000000000000000000000000000000000000000000,
        96'b000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000,
        96'b000000000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000,
        96'b000000000000000000000000001001001001001001001001001000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000001001001001001001001000000000000000000000000000000000000000000000,
        //tile 36, VRAM 54'b000000000000000000000001000011111100111101000000100100
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000001001001001010010010000000000000000000000000000000000000000000000000,
        96'b000000000000000000000001001011100100100100100100100100100100100100000000000000000000000000000000,
        96'b000000000000000000000001001011100100100100100100100100100100100100000000000000000000000000000000,
        96'b000000000000000000001001001011011011011011011011011011011011011011011011011000000000000000000000,
        96'b000000000000000000001001001011011011011011011011011011011011011011011011011000000000000000000000,
        96'b000000000000000000001001001011011011011011011011011011011011011011011011011000000000000000000000,
        96'b000000000000000000001001001001001001001001001001001001000000000000000000000000000000000000000000,
        96'b000000000000001001001001001001001001001001001001001001001000000000000000000000000000000000000000,
        96'b000000000000001001001001001001001001001001001001001001001001000000000000000000000000000000000000,
        96'b000000000000001001001001001001001001001001001001001001001001000000000000000000000000000000000000,
        96'b000000000000000001001001001001001001001001001001001001001001000000000000000000000000000000000000,
        //tile 37, VRAM 54'b000000000000000000000000000001000011111101000000100101
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000001001001010011011011011011011011011011011011011000000000000000000000000000000,
        96'b000000000000000001001001001010011011011011011011011011011011011011000000000000000000000000000000,
        96'b000000000000001001001001001010010010010010010010010010010010010010010010010000000000000000000000,
        96'b000000000000001001001001001010010010010010010010010010010010010010010010010000000000000000000000,
        96'b000000000000001001001001001010010010010010010010010010010010010010010010010000000000000000000000,
        96'b000000001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000,
        96'b000001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000,
        96'b000001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000,
        96'b000001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000,
        96'b000000001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000,
        //tile 38, VRAM 54'b000000000000000000000001000011111100111101000000100110
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000001001001001001001001001001000000000000000000000000000000000000000000000000000000,
        96'b000000000000001001001001001001001001001001001001000000000000000000000000000000000000000000000000,
        96'b000000000001001001001001001001001001001001001001000000000000000000000000000000000000000000000000,
        96'b000000000001001001010001001001001001001001001001001001001000000000000000000000000000000000000000,
        96'b000000000001001001010001001011100100100100100100100100100100100100000000000000000000000000000000,
        96'b000000001001001001010001001011100100100100100100100100100100100100000000000000000000000000000000,
        96'b000001001001001001010010001011011011011011011011011011011011011011011011011000000000000000000000,
        96'b000001001001001001001010001011011011011011011011011011011011011011011011011000000000000000000000,
        96'b000001001001001001001010001011011011011011011011011011011011011011011011011000000000000000000000,
        96'b001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000000,
        96'b001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000,
        96'b001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000,
        96'b001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000,
        96'b001001001001001001001001001001001001001001001001001001001001000000000000000000000000000000000000,
        //tile 39, VRAM 54'b000000000000000000000001000011111100111101000000100111
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000010010001000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000010010010010001000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000010010010001001001001000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000010001001001001001001001010000000000000000000000000000000000000000,
        96'b000000000000000000000000000000010001001001001001001001001000000000000000000000000000000000000000,
        96'b000000000000000000000000000000001001001001001001011100100100100100100100100100100100100000000000,
        96'b000000000000000000000000001001001001001001001001011100100100100100100100100100100100100000000000,
        96'b000000000000000000000000001001001001001001001001011011011011011011011011011011011011011011011011,
        96'b000000000000000000000000001001001001001001001001011011011011011011011011011011011011011011011011,
        96'b000000000000000000000000000000001001001001001001011011011011011011011011011011011011011011011011,
        //tile 40, VRAM 54'b000000000000000000000001000011111100111101000000101000
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000001001001001010010010000000000000000000000000000000000000000000000000,
        96'b000000000000000000000001001001001001001001001001000000000000000000000000000000000000000000000000,
        96'b000000000000000000000001001001001001001001001001000000000000000000000000000000000000000000000000,
        96'b000000000000000000001001001001001010001001001001001000000000000000000000000000000000000000000000,
        96'b000000000000000000001001001010010001001001001001001000000000000000000000000000000000000000000000,
        96'b000000000000000000001001001001001001001001001001001001000000000000000000000000000000000000000000,
        96'b000000000000000000001001001001001001001001001001011100100100100100100100100100100100100000000000,
        96'b000000000000001001001001001001001001001001001001011100100100100100100100100100100100100000000000,
        96'b000000000000001001001001001001001001001001001001011011011011011011011011011011011011011011011011,
        96'b000000000000001001001001001001001001001001001001011011011011011011011011011011011011011011011011,
        96'b000000000000000001001001001001001001001001001001011011011011011011011011011011011011011011011011,
        //tile 41, VRAM 54'b000000000000000000000001000011111100111101000000101001
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000001001001001001000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000001001001001001001001001001001000000000000000000000000000000000000000000000000,
        96'b000000000000000001001001001001001001001001001001000000000000000000000000000000000000000000000000,
        96'b000000000000001001001001001001001001001001001001001000000000000000000000000000000000000000000000,
        96'b000000000000001001001001001001001001001001001001001001010000000000000000000000000000000000000000,
        96'b000000000000001001001001001001001001001001001001001001001000000000000000000000000000000000000000,
        96'b000000001001001001001001001001001001001001001001011100100100100100100100100100100100100000000000,
        96'b000001001001001001001001001001001001001001001001011100100100100100100100100100100100100000000000,
        96'b000001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011,
        96'b000001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011,
        96'b000000001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011,
        //tile 42, VRAM 54'b000000000000000000000001000011111100111101000000101010
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        96'b000000000000000001001001001001001001001001000000000000000000000000000000000000000000000000000000,
        96'b000000000000001001001001001001001001001001001001000000000000000000000000000000000000000000000000,
        96'b000000000001001001001001001001001001001001001001000000000000000000000000000000000000000000000000,
        96'b000000000001001001010001001001001001001001001001001001001000000000000000000000000000000000000000,
        96'b000000000001001001010001001001001001001001001001001001001000000000000000000000000000000000000000,
        96'b000000001001001001010001001001001001001001001001001001001000000000000000000000000000000000000000,
        96'b000001001001001001010010001001001001001001001001001001001000000000000000000000000000000000000000,
        96'b000001001001001001001010001001001001001001001001001001001000000000000000000000000000000000000000,
        96'b000001001001001001001010001001001001001001001001001001001000000000000000000000000000000000000000,
        96'b001001001001001001001001001001001001001001001001011100100100100100100100100100100100100000000000,
        96'b001001001001001001001001001001001001001001001001011100100100100100100100100100100100100000000000,
        96'b001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011,
        96'b001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011,
        96'b001001001001001001001001001001001001001001001001011011011011011011011011011011011011011011011011
    
    };

    always_comb
    begin
        data      = DATA[Tile];
        bitmapIdx = 11'd32 * data[5:0] + PixelY;
        bitmap    = BITMAPS[bitmapIdx];
        color     = bitmap[3*(31-PixelX) +: 3];
        pixel     = data[6*color+6 +: 6];
        Data      = (0 < pixel && pixel < 6) ? pixel + PlayerTwo : pixel;
    end

endmodule
